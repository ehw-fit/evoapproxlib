/***
* This code is a part of EvoApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under The MIT License.
* When used, please cite the following article(s): V. Mrazek, R. Hrbacek, Z. Vasicek and L. Sekanina, "EvoApprox8b: Library of approximate adders and multipliers for circuit design and benchmarking of approximation methods". Design, Automation & Test in Europe Conference & Exhibition (DATE), 2017, Lausanne, 2017, pp. 258-261. doi: 10.23919/DATE.2017.7926993 
* This file contains a circuit from evoapprox8b dataset
***/

// Library = cgp-evoapproxlib
// Circuit = mul8_036.v
// Area   (45) = 497.000000
// Delay  (45) = 1.170000
// Power  (45) = 0.247600
// MAE = 157.316530
// MSE = 40937.375000
// MRE = 4.710000 %
// WCE = 875
// WCRE = 200.000000 %
// EP = 98.500000 %

module mul8_036(A, B, O);
  input [7:0] A;
  input [7:0] B;
  output [15:0] O;
  wire [2031:0] N;

  assign N[0] = A[0];
  assign N[1] = A[0];
  assign N[2] = A[1];
  assign N[3] = A[1];
  assign N[4] = A[2];
  assign N[5] = A[2];
  assign N[6] = A[3];
  assign N[7] = A[3];
  assign N[8] = A[4];
  assign N[9] = A[4];
  assign N[10] = A[5];
  assign N[11] = A[5];
  assign N[12] = A[6];
  assign N[13] = A[6];
  assign N[14] = A[7];
  assign N[15] = A[7];
  assign N[16] = B[0];
  assign N[17] = B[0];
  assign N[18] = B[1];
  assign N[19] = B[1];
  assign N[20] = B[2];
  assign N[21] = B[2];
  assign N[22] = B[3];
  assign N[23] = B[3];
  assign N[24] = B[4];
  assign N[25] = B[4];
  assign N[26] = B[5];
  assign N[27] = B[5];
  assign N[28] = B[6];
  assign N[29] = B[6];
  assign N[30] = B[7];
  assign N[31] = B[7];

  AND2X1 n32(.A(N[18]), .B(N[14]), .Y(N[32]));
  assign N[33] = N[32];
  NOR3X1 n36(.A(N[26]), .B(N[12]), .C(N[14]), .Y(N[36]));
  AND2X1 n38(.A(N[6]), .B(N[24]), .Y(N[38]));
  XOR2X1 n40(.A(N[28]), .B(N[28]), .Y(N[40]));
  assign N[41] = N[40];
  NOR2X1 n42(.A(N[33]), .B(N[32]), .Y(N[42]));
  AND2X1 n46(.A(N[2]), .B(N[16]), .Y(N[46]));
  assign N[47] = N[46];
  XOR2X1 n48(.A(N[18]), .B(N[12]), .Y(N[48]));
  assign N[49] = N[48];
  MUX2X1 n50(.A(N[22]), .B(N[32]), .S(N[18]), .Y(N[50]));
  assign N[51] = N[50];
  NAND2X1 n54(.A(N[49]), .B(N[33]), .Y(N[54]));
  assign N[55] = N[54];
  INVX1 n56(.A(N[33]), .Y(N[56]));
  MUX2X1 n62(.A(N[22]), .B(N[32]), .S(N[55]), .Y(N[62]));
  assign N[63] = N[62];
  NOR2X1 n64(.A(N[41]), .B(N[55]), .Y(N[64]));
  assign N[65] = N[64];
  NOR2X1 n70(.A(N[65]), .B(N[42]), .Y(N[70]));
  NOR2X1 n72(.A(N[49]), .B(N[54]), .Y(N[72]));
  assign N[73] = N[72];
  NAND2X1 n76(.A(N[73]), .B(N[70]), .Y(N[76]));
  assign N[77] = N[76];
  NAND3X1 n86(.A(N[47]), .B(N[24]), .C(N[77]), .Y(N[86]));
  OR2X1 n104(.A(N[73]), .B(N[12]), .Y(N[104]));
  assign N[105] = N[104];
  AND2X1 n106(.A(N[63]), .B(N[56]), .Y(N[106]));
  assign N[107] = N[106];
  INVX1 n116(.A(N[105]), .Y(N[116]));
  AND2X1 n120(.A(N[18]), .B(N[70]), .Y(N[120]));
  assign N[121] = N[120];
  FAX1 n130(.A(N[41]), .B(N[4]), .C(N[30]), .YS(N[130]), .YC(N[131]));
  AND2X1 n134(.A(N[14]), .B(N[16]), .Y(N[134]));
  HAX1 n136(.A(N[73]), .B(N[38]), .YS(N[136]), .YC(N[137]));
  OR2X1 n142(.A(N[41]), .B(N[116]), .Y(N[142]));
  FAX1 n144(.A(N[142]), .B(N[54]), .C(N[51]), .YS(N[144]), .YC(N[145]));
  AND2X1 n164(.A(N[145]), .B(N[131]), .Y(N[164]));
  assign N[165] = N[164];
  AND2X1 n208(.A(N[8]), .B(N[18]), .Y(N[208]));
  assign N[209] = N[208];
  INVX1 n214(.A(N[107]), .Y(N[214]));
  assign N[215] = N[214];
  OAI21X1 n222(.A(N[2]), .B(N[0]), .C(N[26]), .Y(N[222]));
  assign N[223] = N[222];
  BUFX2 n232(.A(N[121]), .Y(N[232]));
  assign N[233] = N[232];
  INVX1 n234(.A(N[223]), .Y(N[234]));
  AND2X1 n238(.A(N[12]), .B(N[18]), .Y(N[238]));
  NOR2X1 n246(.A(N[223]), .B(N[234]), .Y(N[246]));
  NOR2X1 n256(.A(N[73]), .B(N[86]), .Y(N[256]));
  assign N[257] = N[256];
  XNOR2X1 n280(.A(N[137]), .B(N[246]), .Y(N[280]));
  assign N[281] = N[280];
  XNOR2X1 n300(.A(N[281]), .B(N[42]), .Y(N[300]));
  assign N[301] = N[300];
  AND2X1 n342(.A(N[10]), .B(N[20]), .Y(N[342]));
  assign N[343] = N[342];
  AND2X1 n356(.A(N[12]), .B(N[20]), .Y(N[356]));
  AND2X1 n372(.A(N[14]), .B(N[20]), .Y(N[372]));
  AND2X1 n446(.A(N[8]), .B(N[22]), .Y(N[446]));
  AND2X1 n460(.A(N[10]), .B(N[22]), .Y(N[460]));
  AND2X1 n476(.A(N[12]), .B(N[22]), .Y(N[476]));
  OR2X1 n488(.A(N[209]), .B(N[70]), .Y(N[488]));
  assign N[489] = N[488];
  AND2X1 n490(.A(N[14]), .B(N[22]), .Y(N[490]));
  OR2X1 n550(.A(N[215]), .B(N[24]), .Y(N[550]));
  AND2X1 n564(.A(N[8]), .B(N[24]), .Y(N[564]));
  AND2X1 n580(.A(N[10]), .B(N[24]), .Y(N[580]));
  assign N[581] = N[580];
  AND2X1 n594(.A(N[12]), .B(N[24]), .Y(N[594]));
  AND2X1 n608(.A(N[14]), .B(N[24]), .Y(N[608]));
  AND2X1 n654(.A(N[4]), .B(N[26]), .Y(N[654]));
  AND2X1 n668(.A(N[6]), .B(N[26]), .Y(N[668]));
  AND2X1 n682(.A(N[8]), .B(N[26]), .Y(N[682]));
  HAX1 n688(.A(N[105]), .B(N[12]), .YS(N[688]), .YC(N[689]));
  AND2X1 n698(.A(N[10]), .B(N[26]), .Y(N[698]));
  OR2X1 n708(.A(N[33]), .B(N[234]), .Y(N[708]));
  assign N[709] = N[708];
  AND2X1 n712(.A(N[12]), .B(N[26]), .Y(N[712]));
  AND2X1 n728(.A(N[14]), .B(N[26]), .Y(N[728]));
  AND2X1 n772(.A(N[4]), .B(N[28]), .Y(N[772]));
  AND2X1 n786(.A(N[6]), .B(N[28]), .Y(N[786]));
  AND2X1 n802(.A(N[8]), .B(N[28]), .Y(N[802]));
  AND2X1 n816(.A(N[10]), .B(N[28]), .Y(N[816]));
  AND2X1 n832(.A(N[12]), .B(N[28]), .Y(N[832]));
  AND2X1 n846(.A(N[14]), .B(N[28]), .Y(N[846]));
  AND2X1 n876(.A(N[2]), .B(N[30]), .Y(N[876]));
  AND2X1 n890(.A(N[4]), .B(N[30]), .Y(N[890]));
  AND2X1 n906(.A(N[6]), .B(N[30]), .Y(N[906]));
  AND2X1 n920(.A(N[8]), .B(N[30]), .Y(N[920]));
  AND2X1 n934(.A(N[10]), .B(N[30]), .Y(N[934]));
  AND2X1 n950(.A(N[12]), .B(N[30]), .Y(N[950]));
  AND2X1 n964(.A(N[14]), .B(N[30]), .Y(N[964]));
  XOR2X1 n980(.A(N[46]), .B(N[698]), .Y(N[980]));
  assign N[981] = N[980];
  NAND2X1 n1022(.A(N[301]), .B(N[54]), .Y(N[1022]));
  assign N[1023] = N[1022];
  BUFX2 n1054(.A(N[121]), .Y(N[1054]));
  assign N[1055] = N[1054];
  FAX1 n1068(.A(N[134]), .B(N[238]), .C(N[343]), .YS(N[1068]), .YC(N[1069]));
  AND2X1 n1082(.A(N[257]), .B(N[356]), .Y(N[1082]));
  HAX1 n1098(.A(N[65]), .B(N[356]), .YS(N[1098]), .YC(N[1099]));
  INVX1 n1126(.A(N[215]), .Y(N[1126]));
  MUX2X1 n1156(.A(N[446]), .B(N[550]), .S(N[654]), .Y(N[1156]));
  assign N[1157] = N[1156];
  FAX1 n1172(.A(N[460]), .B(N[564]), .C(N[668]), .YS(N[1172]), .YC(N[1173]));
  FAX1 n1186(.A(N[476]), .B(N[580]), .C(N[682]), .YS(N[1186]), .YC(N[1187]));
  FAX1 n1202(.A(N[490]), .B(N[594]), .C(N[698]), .YS(N[1202]), .YC(N[1203]));
  HAX1 n1232(.A(N[608]), .B(N[712]), .YS(N[1232]), .YC(N[1233]));
  HAX1 n1246(.A(N[233]), .B(N[981]), .YS(N[1246]), .YC(N[1247]));
  AND2X1 n1306(.A(N[1054]), .B(N[36]), .Y(N[1306]));
  assign N[1307] = N[1306];
  OR2X1 n1320(.A(N[1068]), .B(N[1055]), .Y(N[1320]));
  assign N[1321] = N[1320];
  FAX1 n1334(.A(N[1098]), .B(N[1069]), .C(N[1172]), .YS(N[1334]), .YC(N[1335]));
  FAX1 n1350(.A(N[372]), .B(N[1082]), .C(N[1186]), .YS(N[1350]), .YC(N[1351]));
  FAX1 n1394(.A(N[1157]), .B(N[772]), .C(N[876]), .YS(N[1394]), .YC(N[1395]));
  FAX1 n1408(.A(N[1173]), .B(N[786]), .C(N[890]), .YS(N[1408]), .YC(N[1409]));
  FAX1 n1424(.A(N[1187]), .B(N[802]), .C(N[906]), .YS(N[1424]), .YC(N[1425]));
  FAX1 n1438(.A(N[1203]), .B(N[816]), .C(N[920]), .YS(N[1438]), .YC(N[1439]));
  FAX1 n1454(.A(N[1233]), .B(N[832]), .C(N[934]), .YS(N[1454]), .YC(N[1455]));
  AND2X1 n1468(.A(N[846]), .B(N[950]), .Y(N[1468]));
  HAX1 n1482(.A(N[846]), .B(N[950]), .YS(N[1482]), .YC(N[1483]));
  BUFX2 n1528(.A(N[489]), .Y(N[1528]));
  assign N[1529] = N[1528];
  AND2X1 n1556(.A(N[581]), .B(N[1307]), .Y(N[1556]));
  assign N[1557] = N[1556];
  FAX1 n1572(.A(N[1334]), .B(N[1321]), .C(N[1394]), .YS(N[1572]), .YC(N[1573]));
  FAX1 n1586(.A(N[1350]), .B(N[1335]), .C(N[1408]), .YS(N[1586]), .YC(N[1587]));
  FAX1 n1602(.A(N[1202]), .B(N[1351]), .C(N[1424]), .YS(N[1602]), .YC(N[1603]));
  AND2X1 n1616(.A(N[1232]), .B(N[1438]), .Y(N[1616]));
  HAX1 n1632(.A(N[1232]), .B(N[1438]), .YS(N[1632]), .YC(N[1633]));
  AND2X1 n1646(.A(N[728]), .B(N[1454]), .Y(N[1646]));
  HAX1 n1660(.A(N[728]), .B(N[1454]), .YS(N[1660]), .YC(N[1661]));
  BUFX2 n1676(.A(N[709]), .Y(N[1676]));
  assign N[1677] = N[1676];
  HAX1 n1690(.A(N[1528]), .B(N[1126]), .YS(N[1690]), .YC(N[1691]));
  OR2X1 n1706(.A(N[165]), .B(N[1529]), .Y(N[1706]));
  XOR2X1 n1734(.A(N[1572]), .B(N[1557]), .Y(N[1734]));
  FAX1 n1750(.A(N[1586]), .B(N[1573]), .C(N[1395]), .YS(N[1750]), .YC(N[1751]));
  FAX1 n1764(.A(N[1602]), .B(N[1587]), .C(N[1409]), .YS(N[1764]), .YC(N[1765]));
  FAX1 n1780(.A(N[1632]), .B(N[1603]), .C(N[1425]), .YS(N[1780]), .YC(N[1781]));
  FAX1 n1794(.A(N[1660]), .B(N[1616]), .C(N[1439]), .YS(N[1794]), .YC(N[1795]));
  FAX1 n1808(.A(N[1482]), .B(N[1646]), .C(N[1455]), .YS(N[1808]), .YC(N[1809]));
  AND2X1 n1824(.A(N[964]), .B(N[1468]), .Y(N[1824]));
  HAX1 n1838(.A(N[964]), .B(N[1468]), .YS(N[1838]), .YC(N[1839]));
  OR2X1 n1854(.A(N[1023]), .B(N[1677]), .Y(N[1854]));
  XOR2X1 n1868(.A(N[1706]), .B(N[1691]), .Y(N[1868]));
  OR2X1 n1898(.A(N[1734]), .B(N[688]), .Y(N[1898]));
  BUFX2 n1912(.A(N[1750]), .Y(N[1912]));
  HAX1 n1928(.A(N[1764]), .B(N[1751]), .YS(N[1928]), .YC(N[1929]));
  FAX1 n1942(.A(N[1780]), .B(N[1765]), .C(N[1929]), .YS(N[1942]), .YC(N[1943]));
  FAX1 n1956(.A(N[1794]), .B(N[1781]), .C(N[1943]), .YS(N[1956]), .YC(N[1957]));
  FAX1 n1972(.A(N[1808]), .B(N[1795]), .C(N[1957]), .YS(N[1972]), .YC(N[1973]));
  FAX1 n1986(.A(N[1838]), .B(N[1809]), .C(N[1973]), .YS(N[1986]), .YC(N[1987]));
  OR2X1 n2016(.A(N[1824]), .B(N[1987]), .Y(N[2016]));

  assign O[0] = N[32];
  assign O[1] = N[980];
  assign O[2] = N[1246];
  assign O[3] = N[816];
  assign O[4] = N[1676];
  assign O[5] = N[1854];
  assign O[6] = N[1868];
  assign O[7] = N[1780];
  assign O[8] = N[1898];
  assign O[9] = N[1912];
  assign O[10] = N[1928];
  assign O[11] = N[1942];
  assign O[12] = N[1956];
  assign O[13] = N[1972];
  assign O[14] = N[1986];
  assign O[15] = N[2016];

endmodule



// internal reference: cgp-evoapproxlib.08.mul8_036

