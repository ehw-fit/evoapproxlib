/***
* This code is a part of ApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under a XXXX public license.
* When used, please cite the following article: tbd 
* This file is pareto optimal sub-set in the pdk45_pwr and mae% parameters
***/

module mul12u_pwr_0_146_mae_00_4500(A, B, O);
  input [11:0] A, B;
  output [23:0] O;
  wire n_1418, n_1365, n_458, n_703, n_1385, n_785, n_1049, n_787, n_43, n_1043;
  wire n_789, n_1045, n_1047, n_1287, n_1285, n_1283, n_1281, n_145, n_1289, n_1502;
  wire n_1518, n_889, n_1248, n_1443, n_1051, n_1391, n_1357, n_1180, n_1352, n_1182;
  wire n_1496, n_949, n_1508, n_39, n_1395, n_393, n_1467, n_1397, n_1512, n_1510;
  wire n_1516, n_1514, n_1022, n_1457, n_433, n_1020, n_1027, n_1024, n_1025, n_1379;
  wire n_23, n_22, n_21, n_20, n_27, n_26, n_24, n_8, n_29, n_28;
  wire n_1225, n_1377, n_1260, n_1465, n_1156, n_891, n_1400, n_893, n_1414, n_895;
  wire n_894, n_897, n_658, n_656, n_1408, n_1030, n_1270, n_1141, n_1231, n_635;
  wire n_1277, n_1402, n_1404, n_633, n_1481, n_934, n_1484, n_1275, n_18, n_19;
  wire n_16, n_17, n_14, n_15, n_12, n_13, n_10, n_11, n_96, n_1482;
  wire n_98, n_883, n_881, n_887, n_527, n_885, n_137, n_643, n_1242, n_357;
  wire n_1008, n_1129, n_1004, n_1006, n_1000, n_1305, n_1002, n_1488, n_1158, n_1498;
  wire n_1152, n_1268, n_1150, n_1494, n_1143, n_1492, n_1154, n_1490, n_81, n_80;
  wire n_85, n_1123, n_734, n_1504, n_1522, n_1520, n_107, n_1250, n_1018, n_1254;
  wire n_1256, n_1012, n_1010, n_1016, n_615, n_1014, n_1149, n_918, n_1309, n_852;
  wire n_914, n_1311, n_916, n_1313, n_1145, n_1500, n_1147, n_115, n_1393, n_78;
  wire n_79, n_1131, n_1399, n_1506, n_217, n_1416, n_1133, n_213, n_1412, n_1410;
  wire n_503, n_219, n_920, n_275, n_274, n_1176, n_1304, n_271, n_1301, n_1264;
  wire n_1406, n_1266, n_1137, n_1178, n_371, n_1262, n_1486, n_1252, n_1139, n_1174;
  wire n_165, n_167, n_649, n_1387, n_65, n_1383, n_1381, n_1463, n_1307, n_756;
  wire n_1451, n_1258, n_1303, n_209, n_758, n_1469, n_1373, n_1279, n_1371, n_262;
  wire n_9, n_1375, n_4, n_5, n_6, n_7, n_0, n_1, n_2, n_3;
  wire n_1135, n_1272, n_1420, n_879, n_59, n_1389, n_174, n_178, n_51, n_1274;
  wire n_1471, n_1473, n_1475, n_1477, n_1479, n_766, n_764, n_762, n_760;
  assign n_0 = A[0];
  assign n_1 = A[1];
  assign n_2 = A[2];
  assign n_3 = A[3];
  assign n_4 = A[4];
  assign n_5 = A[5];
  assign n_6 = A[6];
  assign n_7 = A[7];
  assign n_8 = A[8];
  assign n_9 = A[9];
  assign n_10 = A[10];
  assign n_11 = A[11];
  assign n_12 = B[0];
  assign n_13 = B[1];
  assign n_14 = B[2];
  assign n_15 = B[3];
  assign n_16 = B[4];
  assign n_17 = B[5];
  assign n_18 = B[6];
  assign n_19 = B[7];
  assign n_20 = B[8];
  assign n_21 = B[9];
  assign n_22 = B[10];
  assign n_23 = B[11];
  assign n_24 = n_13 & n_22;
  assign n_26 = n_7 & n_24;
  assign n_27 = n_23 & n_26;
  assign n_28 = n_18 ^ n_18;
  assign n_29 = n_5 & n_27;
  assign n_39 = ~n_28;
  assign n_43 = n_5 & n_27;
  assign n_51 = n_43;
  assign n_59 = n_28;
  assign n_65 = n_28 & n_13;
  assign n_78 = n_29 ^ n_51;
  assign n_79 = n_39;
  assign n_80 = n_1 & n_78;
  assign n_81 = n_6 & n_9;
  assign n_85 = n_5 & n_80;
  assign n_96 = n_13 & n_78;
  assign n_98 = ~(n_79 | n_6);
  assign n_107 = ~n_85;
  assign n_115 = n_17 & n_85;
  assign n_137 = n_96 & n_14;
  assign n_145 = n_22 & n_78;
  assign n_165 = n_78 & n_78;
  assign n_167 = ~n_165;
  assign n_174 = ~n_145;
  assign n_178 = ~n_65;
  assign n_209 = ~(n_10 | n_167);
  assign n_213 = n_81 & n_22;
  assign n_217 = ~(n_65 | n_78);
  assign n_219 = n_98;
  assign n_262 = ~(n_9 & n_80);
  assign n_271 = ~n_39;
  assign n_274 = ~n_271;
  assign n_275 = ~n_137;
  assign n_357 = ~(n_107 | n_262);
  assign n_371 = ~n_145;
  assign n_393 = n_219 & n_165;
  assign n_433 = ~(n_275 | n_3);
  assign n_458 = ~n_59;
  assign n_503 = ~n_262;
  assign n_527 = n_11 & n_17;
  assign n_615 = ~n_458;
  assign n_633 = ~(n_219 | n_219);
  assign n_635 = n_271;
  assign n_643 = n_98;
  assign n_649 = n_643 & n_7;
  assign n_656 = n_10 & n_18;
  assign n_658 = n_11 & n_18;
  assign n_703 = ~n_137;
  assign n_734 = ~n_615;
  assign n_756 = n_213;
  assign n_758 = ~n_635;
  assign n_760 = n_527 & n_656;
  assign n_762 = n_393 & n_635;
  assign n_764 = n_758 | n_174;
  assign n_766 = n_760 | n_762;
  assign n_785 = n_9 & n_213;
  assign n_787 = n_10 & n_19;
  assign n_789 = n_11 & n_19;
  assign n_852 = n_209 & n_178;
  assign n_879 = ~(n_764 & n_785);
  assign n_881 = n_764 & n_785;
  assign n_883 = n_879 & n_756;
  assign n_885 = n_879 ^ n_756;
  assign n_887 = n_881 | n_883;
  assign n_889 = n_658 ^ n_787;
  assign n_891 = n_658 & n_787;
  assign n_893 = n_889 & n_766;
  assign n_894 = ~n_217;
  assign n_895 = n_889 ^ n_766;
  assign n_897 = n_891 | n_893;
  assign n_914 = n_8 & n_20;
  assign n_916 = n_9 & n_20;
  assign n_918 = n_10 & n_20;
  assign n_920 = n_11 & n_20;
  assign n_934 = ~n_85;
  assign n_949 = n_145 & n_633;
  assign n_1000 = n_949;
  assign n_1002 = n_885 & n_914;
  assign n_1004 = n_1000;
  assign n_1006 = ~n_1000;
  assign n_1008 = n_1002;
  assign n_1010 = n_895 ^ n_916;
  assign n_1012 = n_895 & n_916;
  assign n_1014 = n_1010 & n_887;
  assign n_1016 = n_1010 ^ n_887;
  assign n_1018 = n_1012 | n_1014;
  assign n_1020 = n_789 ^ n_918;
  assign n_1022 = n_789 & n_918;
  assign n_1024 = n_1020 & n_897;
  assign n_1025 = n_1020 ^ n_897;
  assign n_1027 = n_1022 ^ n_1024;
  assign n_1030 = ~n_371;
  assign n_1043 = n_7 & n_21;
  assign n_1045 = n_8 & n_21;
  assign n_1047 = n_9 & n_21;
  assign n_1049 = n_10 & n_21;
  assign n_1051 = n_11 & n_21;
  assign n_1123 = n_1006 & n_1043;
  assign n_1129 = n_1123 | n_96;
  assign n_1131 = n_1016 ^ n_1045;
  assign n_1133 = n_1016 & n_1045;
  assign n_1135 = n_1131 & n_1008;
  assign n_1137 = n_1131 ^ n_1008;
  assign n_1139 = n_1133 | n_1135;
  assign n_1141 = n_1025 ^ n_1047;
  assign n_1143 = n_1025 & n_1047;
  assign n_1145 = n_1141 & n_1018;
  assign n_1147 = n_1141 ^ n_1018;
  assign n_1149 = n_1143 | n_1145;
  assign n_1150 = n_920 ^ n_1049;
  assign n_1152 = n_920 & n_1049;
  assign n_1154 = n_1150 & n_1027;
  assign n_1156 = n_1150 ^ n_1027;
  assign n_1158 = n_1152 | n_1154;
  assign n_1174 = n_7 & n_22;
  assign n_1176 = n_8 & n_22;
  assign n_1178 = n_9 & n_22;
  assign n_1180 = n_10 & n_22;
  assign n_1182 = n_11 & n_22;
  assign n_1225 = ~(n_1006 | n_1030);
  assign n_1231 = ~n_1225;
  assign n_1242 = ~n_165;
  assign n_1248 = n_1242;
  assign n_1250 = ~n_209;
  assign n_1252 = n_1137 ^ n_1174;
  assign n_1254 = n_1137 & n_1174;
  assign n_1256 = n_1252 & n_1129;
  assign n_1258 = n_1252 ^ n_1129;
  assign n_1260 = n_1254 | n_1256;
  assign n_1262 = n_1147 ^ n_1176;
  assign n_1264 = n_1147 & n_1176;
  assign n_1266 = n_1262 & n_1139;
  assign n_1268 = n_1262 ^ n_1139;
  assign n_1270 = n_1264 | n_1266;
  assign n_1272 = n_1156 ^ n_1178;
  assign n_1274 = n_1156 & n_1178;
  assign n_1275 = n_1272 & n_1149;
  assign n_1277 = n_1272 ^ n_1149;
  assign n_1279 = n_1274 ^ n_1275;
  assign n_1281 = n_1051 ^ n_1180;
  assign n_1283 = n_1051 & n_1180;
  assign n_1285 = n_1281 & n_1158;
  assign n_1287 = n_1281 ^ n_1158;
  assign n_1289 = n_1283 | n_1285;
  assign n_1301 = n_5 & n_23;
  assign n_1303 = n_6 & n_23;
  assign n_1304 = n_357;
  assign n_1305 = n_7 & n_23;
  assign n_1307 = n_8 & n_23;
  assign n_1309 = n_9 & n_23;
  assign n_1311 = n_10 & n_23;
  assign n_1313 = n_11 & n_23;
  assign n_1352 = n_21 | n_274;
  assign n_1357 = ~(n_1030 | n_1231);
  assign n_1365 = n_1248 & n_1301;
  assign n_1371 = n_1365;
  assign n_1373 = n_1258 ^ n_1303;
  assign n_1375 = n_1258;
  assign n_1377 = n_1373 & n_458;
  assign n_1379 = ~(n_1373 & n_1250);
  assign n_1381 = n_1375 | n_1377;
  assign n_1383 = n_1268 ^ n_1305;
  assign n_1385 = n_1268 & n_1305;
  assign n_1387 = n_1383 & n_1260;
  assign n_1389 = n_1383 ^ n_1260;
  assign n_1391 = n_1385 ^ n_1387;
  assign n_1393 = n_1277 ^ n_1307;
  assign n_1395 = n_1277 & n_1307;
  assign n_1397 = n_1393 & n_1270;
  assign n_1399 = n_1393 ^ n_1270;
  assign n_1400 = n_1395 | n_1397;
  assign n_1402 = n_1287 ^ n_1309;
  assign n_1404 = n_1287 & n_1309;
  assign n_1406 = n_1402 & n_1279;
  assign n_1408 = n_1402 ^ n_1279;
  assign n_1410 = n_1404 | n_1406;
  assign n_1412 = n_1182 ^ n_1311;
  assign n_1414 = n_1182 & n_1311;
  assign n_1416 = n_1412 & n_1289;
  assign n_1418 = n_1412 ^ n_1289;
  assign n_1420 = n_1414 | n_1416;
  assign n_1443 = ~n_78;
  assign n_1451 = ~(n_934 & n_1443);
  assign n_1457 = ~(n_1352 | n_649);
  assign n_1463 = n_1457;
  assign n_1465 = n_1379 ^ n_1371;
  assign n_1467 = n_1379 & n_1371;
  assign n_1469 = n_174 & n_1463;
  assign n_1471 = n_1465;
  assign n_1473 = n_1467 | n_1469;
  assign n_1475 = n_1389 ^ n_1381;
  assign n_1477 = n_1389 & n_1381;
  assign n_1479 = n_1475 & n_1473;
  assign n_1481 = n_1475 ^ n_1473;
  assign n_1482 = n_1477 | n_1479;
  assign n_1484 = n_1399 ^ n_1391;
  assign n_1486 = n_1399 & n_1391;
  assign n_1488 = n_1484 & n_1482;
  assign n_1490 = n_1484 ^ n_1482;
  assign n_1492 = n_1486 | n_1488;
  assign n_1494 = n_1408 ^ n_1400;
  assign n_1496 = n_1408 & n_1400;
  assign n_1498 = n_1494 & n_1492;
  assign n_1500 = n_1494 ^ n_1492;
  assign n_1502 = n_1496 | n_1498;
  assign n_1504 = n_1418 ^ n_1410;
  assign n_1506 = n_1418 & n_1410;
  assign n_1508 = n_1504 & n_1502;
  assign n_1510 = n_1504 ^ n_1502;
  assign n_1512 = n_1506 | n_1508;
  assign n_1514 = n_1313 ^ n_1420;
  assign n_1516 = n_1313 & n_1420;
  assign n_1518 = n_1514 & n_1512;
  assign n_1520 = n_1514 ^ n_1512;
  assign n_1522 = n_1516 | n_1518;
  assign O[0] = n_1357;
  assign O[1] = n_894;
  assign O[2] = n_115;
  assign O[3] = n_1304;
  assign O[4] = n_1;
  assign O[5] = n_98;
  assign O[6] = n_703;
  assign O[7] = n_1004;
  assign O[8] = n_357;
  assign O[9] = n_1418;
  assign O[10] = n_503;
  assign O[11] = n_852;
  assign O[12] = n_1469;
  assign O[13] = n_734;
  assign O[14] = n_107;
  assign O[15] = n_1451;
  assign O[16] = n_433;
  assign O[17] = n_1471;
  assign O[18] = n_1481;
  assign O[19] = n_1490;
  assign O[20] = n_1500;
  assign O[21] = n_1510;
  assign O[22] = n_1520;
  assign O[23] = n_1522;
endmodule


// internal reference: cgp-compare17.12.mul12u_pwr_0_146_mae_00_4500

