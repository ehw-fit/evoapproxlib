/***
    * This code is a part of ApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under a XXXX public license.
    * When used, please cite the following article: tbd 
    * This file is pareto optimal sub-set in the pwr and mae parameters
    ***/
    
// ../../../cgp.nn/res/11b_160129\rcam\e01.0\run.00093.txt
module mul11u_pwr_0_367_mae_00_2508(A, B, O);
  input [10:0] A, B;
  output [21:0] O;
  wire [10:0] A, B;
  wire [21:0] O;
  wire sig_33, sig_103, sig_152, sig_155, sig_166, sig_210;
  wire sig_213, sig_214, sig_215, sig_216, sig_217, sig_218;
  wire sig_227, sig_228, sig_229, sig_268, sig_270, sig_271;
  wire sig_272, sig_273, sig_274, sig_275, sig_277, sig_278;
  wire sig_279, sig_280, sig_281, sig_289, sig_290, sig_291;
  wire sig_292, sig_322, sig_325, sig_326, sig_328, sig_329;
  wire sig_330, sig_331, sig_332, sig_333, sig_334, sig_335;
  wire sig_336, sig_337, sig_338, sig_339, sig_340, sig_341;
  wire sig_342, sig_343, sig_344, sig_351, sig_352, sig_354;
  wire sig_355, sig_381, sig_383, sig_384, sig_385, sig_386;
  wire sig_387, sig_388, sig_389, sig_390, sig_391, sig_392;
  wire sig_393, sig_394, sig_395, sig_396, sig_397, sig_398;
  wire sig_399, sig_401, sig_402, sig_403, sig_404, sig_406;
  wire sig_407, sig_414, sig_416, sig_417, sig_418, sig_437;
  wire sig_440, sig_441, sig_442, sig_443, sig_444, sig_445;
  wire sig_446, sig_447, sig_448, sig_449, sig_450, sig_451;
  wire sig_452, sig_453, sig_454, sig_455, sig_456, sig_457;
  wire sig_458, sig_459, sig_460, sig_461, sig_462, sig_463;
  wire sig_464, sig_465, sig_466, sig_467, sig_469, sig_470;
  wire sig_474, sig_475, sig_476, sig_477, sig_478, sig_479;
  wire sig_480, sig_481, sig_495, sig_498, sig_499, sig_500;
  wire sig_501, sig_502, sig_503, sig_504, sig_505, sig_506;
  wire sig_507, sig_508, sig_509, sig_510, sig_511, sig_512;
  wire sig_513, sig_514, sig_515, sig_516, sig_517, sig_518;
  wire sig_519, sig_520, sig_521, sig_522, sig_523, sig_524;
  wire sig_525, sig_526, sig_527, sig_529, sig_530, sig_531;
  wire sig_532, sig_533, sig_536, sig_537, sig_538, sig_539;
  wire sig_540, sig_541, sig_542, sig_543, sig_544, sig_551;
  wire sig_552, sig_553, sig_554, sig_556, sig_557, sig_558;
  wire sig_559, sig_560, sig_561, sig_562, sig_563, sig_564;
  wire sig_565, sig_566, sig_567, sig_568, sig_569, sig_570;
  wire sig_571, sig_572, sig_573, sig_574, sig_575, sig_576;
  wire sig_577, sig_578, sig_579, sig_580, sig_581, sig_583;
  wire sig_584, sig_585, sig_586, sig_587, sig_588, sig_589;
  wire sig_590, sig_591, sig_592, sig_593, sig_594, sig_595;
  wire sig_596, sig_598, sig_599, sig_600, sig_601, sig_602;
  wire sig_603, sig_604, sig_605, sig_606, sig_607, sig_611;
  wire sig_614, sig_615, sig_616, sig_617, sig_619, sig_620;
  wire sig_621, sig_622, sig_624, sig_625, sig_626, sig_627;
  wire sig_629, sig_630, sig_631, sig_632, sig_634, sig_635;
  wire sig_636, sig_637, sig_639, sig_640, sig_641, sig_642;
  wire sig_644, sig_645, sig_646, sig_647, sig_649, sig_650;
  wire sig_651, sig_652, sig_654, sig_655, sig_656, sig_657;
  assign sig_33 = A[0] & B[1];
  assign O[1] = A[0] & sig_33;
  assign sig_103 = A[10];
  assign sig_152 = B[3] & sig_103;
  assign sig_155 = sig_152 & B[2];
  assign sig_166 = A[10] & B[3];
  assign sig_210 = A[9] & B[4];
  assign sig_213 = sig_210;
  assign sig_214 = sig_155 ^ sig_166;
  assign sig_215 = sig_155;
  assign sig_216 = sig_214 & sig_213;
  assign sig_217 = sig_214 ^ sig_213;
  assign sig_218 = sig_215 | sig_216;
  assign sig_227 = A[8] & B[8];
  assign sig_228 = A[9] & B[4];
  assign sig_229 = A[10] & B[4];
  assign sig_268 = A[9] & sig_227;
  assign sig_270 = B[2] & A[10];
  assign sig_271 = sig_268;
  assign sig_272 = sig_217 ^ sig_228;
  assign sig_273 = sig_217 & sig_228;
  assign sig_274 = sig_272 & sig_271;
  assign sig_275 = sig_272 ^ sig_271;
  assign O[6] = sig_273 | sig_274;
  assign sig_277 = sig_218 ^ sig_229;
  assign sig_278 = sig_218 & sig_229;
  assign sig_279 = sig_277 & O[6];
  assign sig_280 = sig_277 ^ O[6];
  assign sig_281 = sig_278 | sig_279;
  assign sig_289 = A[7] & B[5];
  assign sig_290 = A[8] & B[5];
  assign sig_291 = A[9] & B[5];
  assign sig_292 = A[10] & B[5];
  assign sig_322 = A[3] & A[3];
  assign O[5] = B[2] & sig_322;
  assign sig_325 = sig_270 | sig_289;
  assign sig_326 = B[7] & sig_289;
  assign sig_328 = sig_325 ^ O[5];
  assign sig_329 = sig_326;
  assign sig_330 = sig_275 ^ sig_290;
  assign sig_331 = sig_275 & sig_290;
  assign sig_332 = sig_330 & sig_329;
  assign sig_333 = sig_330 ^ sig_329;
  assign sig_334 = sig_331 | sig_332;
  assign sig_335 = sig_280 ^ sig_291;
  assign sig_336 = sig_280 & sig_291;
  assign sig_337 = sig_335 & sig_334;
  assign sig_338 = sig_335 ^ sig_334;
  assign sig_339 = sig_336 | sig_337;
  assign sig_340 = sig_281 ^ sig_292;
  assign sig_341 = sig_281 & sig_292;
  assign sig_342 = sig_340 & sig_339;
  assign sig_343 = sig_340 ^ sig_339;
  assign sig_344 = sig_341 | sig_342;
  assign sig_351 = A[6] & B[6];
  assign sig_352 = A[7] & B[6];
  assign O[11] = A[8] & B[6];
  assign sig_354 = A[9] & B[6];
  assign sig_355 = A[10] & B[6];
  assign sig_381 = B[5] & A[10];
  assign sig_383 = sig_328 ^ sig_351;
  assign sig_384 = B[0] & sig_351;
  assign sig_385 = A[5] & B[2];
  assign sig_386 = sig_383;
  assign sig_387 = sig_384 | sig_385;
  assign sig_388 = sig_333 ^ sig_352;
  assign sig_389 = sig_333 & sig_352;
  assign sig_390 = sig_388 & sig_387;
  assign sig_391 = sig_388 ^ sig_387;
  assign sig_392 = sig_389 | sig_390;
  assign sig_393 = sig_338 ^ O[11];
  assign sig_394 = sig_338 & O[11];
  assign sig_395 = sig_393 & sig_392;
  assign sig_396 = sig_393 ^ sig_392;
  assign sig_397 = sig_394 | sig_395;
  assign sig_398 = sig_343 ^ sig_354;
  assign sig_399 = sig_343 & sig_354;
  assign O[8] = sig_398 & sig_397;
  assign sig_401 = sig_398 ^ sig_397;
  assign sig_402 = sig_399 | O[8];
  assign sig_403 = sig_344 ^ sig_355;
  assign sig_404 = sig_344 & sig_355;
  assign O[9] = sig_403 & sig_402;
  assign sig_406 = sig_403 ^ sig_402;
  assign sig_407 = sig_404 | O[9];
  assign sig_414 = A[6] & B[7];
  assign O[3] = A[7] & B[7];
  assign sig_416 = A[8] & B[7];
  assign sig_417 = A[9] & B[7];
  assign sig_418 = A[10] & B[7];
  assign sig_437 = sig_381 & A[8];
  assign sig_440 = sig_437;
  assign sig_441 = sig_386;
  assign sig_442 = B[7] & A[6];
  assign sig_443 = sig_441 ^ sig_440;
  assign sig_444 = sig_441 ^ sig_440;
  assign sig_445 = sig_442 | sig_443;
  assign sig_446 = sig_391 | sig_414;
  assign sig_447 = sig_391 | sig_414;
  assign sig_448 = sig_446 & B[6];
  assign sig_449 = sig_446 ^ sig_445;
  assign sig_450 = sig_447 | sig_448;
  assign sig_451 = sig_396 ^ O[3];
  assign sig_452 = sig_396 & O[3];
  assign sig_453 = sig_451 & sig_450;
  assign sig_454 = sig_451 ^ sig_450;
  assign sig_455 = sig_452 | sig_453;
  assign sig_456 = sig_401 ^ sig_416;
  assign sig_457 = sig_401 & sig_416;
  assign sig_458 = sig_456 & sig_455;
  assign sig_459 = sig_456 ^ sig_455;
  assign sig_460 = sig_457 | sig_458;
  assign sig_461 = sig_406 ^ sig_417;
  assign sig_462 = sig_406 & sig_417;
  assign sig_463 = sig_461 & sig_460;
  assign sig_464 = sig_461 ^ sig_460;
  assign sig_465 = sig_462 | sig_463;
  assign sig_466 = sig_407 ^ sig_418;
  assign sig_467 = sig_407 & sig_418;
  assign O[0] = sig_466 & sig_465;
  assign sig_469 = sig_466 ^ sig_465;
  assign sig_470 = sig_467 | O[0];
  assign sig_474 = A[8] & B[8];
  assign sig_475 = A[4] & B[8];
  assign sig_476 = A[5] & B[8];
  assign sig_477 = A[6] & B[8];
  assign sig_478 = A[7] & B[8];
  assign sig_479 = A[8] & B[8];
  assign sig_480 = A[9] & B[8];
  assign sig_481 = A[10] & B[8];
  assign sig_495 = B[7] & sig_474;
  assign sig_498 = sig_495;
  assign sig_499 = sig_444 | sig_475;
  assign sig_500 = sig_444;
  assign sig_501 = sig_499 & sig_498;
  assign sig_502 = sig_499 ^ sig_498;
  assign sig_503 = sig_500 | sig_501;
  assign sig_504 = sig_449 ^ sig_476;
  assign sig_505 = sig_449 & sig_476;
  assign sig_506 = sig_504 & sig_503;
  assign sig_507 = sig_504 ^ sig_503;
  assign sig_508 = sig_505 | sig_506;
  assign sig_509 = sig_454 ^ sig_477;
  assign sig_510 = sig_454 & sig_477;
  assign sig_511 = sig_509 & sig_508;
  assign sig_512 = sig_509 ^ sig_508;
  assign sig_513 = sig_510 ^ sig_511;
  assign sig_514 = sig_459 ^ sig_478;
  assign sig_515 = sig_459 & sig_478;
  assign sig_516 = sig_514 & sig_513;
  assign sig_517 = sig_514 ^ sig_513;
  assign sig_518 = sig_515 | sig_516;
  assign sig_519 = sig_464 ^ sig_479;
  assign sig_520 = sig_464 & sig_479;
  assign sig_521 = sig_519 & sig_518;
  assign sig_522 = sig_519 ^ sig_518;
  assign sig_523 = sig_520 ^ sig_521;
  assign sig_524 = sig_469 ^ sig_480;
  assign sig_525 = sig_469 & sig_480;
  assign sig_526 = sig_524 & sig_523;
  assign sig_527 = sig_524 ^ sig_523;
  assign O[2] = sig_525 ^ sig_526;
  assign sig_529 = sig_470 ^ sig_481;
  assign sig_530 = sig_470 & sig_481;
  assign sig_531 = sig_529 & O[2];
  assign sig_532 = sig_529 ^ O[2];
  assign sig_533 = sig_530 | sig_531;
  assign sig_536 = A[9] & B[8];
  assign sig_537 = A[3] & B[9];
  assign sig_538 = A[4] & B[9];
  assign sig_539 = A[5] & B[9];
  assign sig_540 = A[6] & B[9];
  assign sig_541 = A[7] & B[9];
  assign sig_542 = A[8] & B[9];
  assign sig_543 = A[9] & B[9];
  assign sig_544 = A[10] & B[9];
  assign sig_551 = A[5];
  assign sig_552 = B[3] ^ sig_536;
  assign sig_553 = B[4] & A[1];
  assign sig_554 = sig_552 & sig_551;
  assign sig_556 = sig_553 | sig_554;
  assign sig_557 = sig_502 ^ sig_537;
  assign sig_558 = sig_502 & sig_537;
  assign sig_559 = sig_557 & sig_556;
  assign sig_560 = sig_557 ^ sig_556;
  assign sig_561 = sig_558 | sig_559;
  assign sig_562 = sig_507 ^ sig_538;
  assign sig_563 = sig_507 & sig_538;
  assign sig_564 = sig_562 & sig_561;
  assign sig_565 = sig_562 ^ sig_561;
  assign sig_566 = sig_563 | sig_564;
  assign sig_567 = sig_512 ^ sig_539;
  assign sig_568 = sig_512 & sig_539;
  assign sig_569 = sig_567 & sig_566;
  assign sig_570 = sig_567 ^ sig_566;
  assign sig_571 = sig_568 | sig_569;
  assign sig_572 = sig_517 ^ sig_540;
  assign sig_573 = sig_517 & sig_540;
  assign sig_574 = sig_572 & sig_571;
  assign sig_575 = sig_572 ^ sig_571;
  assign sig_576 = sig_573 | sig_574;
  assign sig_577 = sig_522 ^ sig_541;
  assign sig_578 = sig_522 & sig_541;
  assign sig_579 = sig_577 & sig_576;
  assign sig_580 = sig_577 ^ sig_576;
  assign sig_581 = sig_578 | sig_579;
  assign O[10] = sig_527 ^ sig_542;
  assign sig_583 = sig_527 & sig_542;
  assign sig_584 = O[10] & sig_581;
  assign sig_585 = O[10] ^ sig_581;
  assign sig_586 = sig_583 | sig_584;
  assign sig_587 = sig_532 ^ sig_543;
  assign sig_588 = sig_532 & sig_543;
  assign sig_589 = sig_587 & sig_586;
  assign sig_590 = sig_587 ^ sig_586;
  assign sig_591 = sig_588 | sig_589;
  assign sig_592 = sig_533 ^ sig_544;
  assign sig_593 = sig_533 & sig_544;
  assign sig_594 = sig_592 & sig_591;
  assign sig_595 = sig_592 ^ sig_591;
  assign sig_596 = sig_593 | sig_594;
  assign sig_598 = A[9] & A[2];
  assign sig_599 = A[2] & B[10];
  assign sig_600 = A[3] & B[10];
  assign sig_601 = A[4] & B[10];
  assign sig_602 = A[5] & B[10];
  assign sig_603 = A[6] & B[10];
  assign sig_604 = A[7] & B[10];
  assign sig_605 = A[8] & B[10];
  assign sig_606 = A[9] & B[10];
  assign sig_607 = A[10] & B[10];
  assign sig_611 = B[7] & sig_598;
  assign sig_614 = sig_611;
  assign sig_615 = sig_560 ^ sig_599;
  assign sig_616 = sig_560 & sig_599;
  assign sig_617 = sig_615 & sig_614;
  assign O[12] = sig_615 ^ sig_614;
  assign sig_619 = sig_616 ^ sig_617;
  assign sig_620 = sig_565 ^ sig_600;
  assign sig_621 = sig_565 & sig_600;
  assign sig_622 = sig_620 & sig_619;
  assign O[13] = sig_620 ^ sig_619;
  assign sig_624 = sig_621 ^ sig_622;
  assign sig_625 = sig_570 ^ sig_601;
  assign sig_626 = sig_570 & sig_601;
  assign sig_627 = sig_625 & sig_624;
  assign O[14] = sig_625 ^ sig_624;
  assign sig_629 = sig_626 | sig_627;
  assign sig_630 = sig_575 ^ sig_602;
  assign sig_631 = sig_575 & sig_602;
  assign sig_632 = sig_630 & sig_629;
  assign O[15] = sig_630 ^ sig_629;
  assign sig_634 = sig_631 | sig_632;
  assign sig_635 = sig_580 ^ sig_603;
  assign sig_636 = sig_580 & sig_603;
  assign sig_637 = sig_635 & sig_634;
  assign O[4] = sig_635 ^ sig_634;
  assign sig_639 = sig_636 | sig_637;
  assign sig_640 = sig_585 ^ sig_604;
  assign sig_641 = sig_585 & sig_604;
  assign sig_642 = sig_640 & sig_639;
  assign O[17] = sig_640 ^ sig_639;
  assign sig_644 = sig_641 ^ sig_642;
  assign sig_645 = sig_590 ^ sig_605;
  assign sig_646 = sig_590 & sig_605;
  assign sig_647 = sig_645 & sig_644;
  assign O[18] = sig_645 ^ sig_644;
  assign sig_649 = sig_646 | sig_647;
  assign sig_650 = sig_595 ^ sig_606;
  assign sig_651 = sig_595 & sig_606;
  assign sig_652 = sig_650 & sig_649;
  assign O[19] = sig_650 ^ sig_649;
  assign sig_654 = sig_651 | sig_652;
  assign sig_655 = sig_596 ^ sig_607;
  assign sig_656 = sig_596 & sig_607;
  assign sig_657 = sig_655 & sig_654;
  assign O[20] = sig_655 ^ sig_654;
  assign O[21] = sig_656 | sig_657;
  assign O[7] = O[3]; // default output
  assign O[16] = O[4]; // default output
endmodule


// internal reference: cgp-nn-iccad16.11.mul11u_pwr_0_367_mae_00_2508

