/***
* This code is a part of EvoApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under The MIT License.
* When used, please cite the following article(s): Z. Vasicek and L. Sekanina, "Evolutionary Approach to Approximate Digital Circuits Design" in IEEE Transactions on Evolutionary Computation, vol. 19, no. 3, pp. 432-444, June 2015. doi: 10.1109/TEVC.2014.2336175 
* This file contains a circuit from a sub-set of pareto optimal circuits with respect to the pwr and ep parameters
***/
// MAE% = 1.39 %
// MAE = 59650503 
// WCE% = 22.22 %
// WCE = 954408050 
// WCRE% = 22.22 %
// EP% = 80.98 %
// MRE% = 3.32 %
// MSE = 27897.246e12 
// PDK45_PWR = 1.984 mW
// PDK45_AREA = 3094.1 um2
// PDK45_DELAY = 3.23 ns

module mul16u_0Z6 (
    A,
    B,
    O
);

input [15:0] A;
input [15:0] B;
output [31:0] O;

wire sig_32,sig_33,sig_34,sig_35,sig_36,sig_37,sig_38,sig_39,sig_40,sig_41,sig_42,sig_43,sig_44,sig_45,sig_46,sig_47,sig_48,sig_49,sig_50,sig_51;
wire sig_56,sig_58,sig_63,sig_65,sig_66,sig_67,sig_69,sig_71,sig_75,sig_80,sig_82,sig_83,sig_85,sig_98,sig_100,sig_102,sig_104,sig_105,sig_106,sig_107;
wire sig_108,sig_109,sig_111,sig_113,sig_117,sig_122,sig_123,sig_124,sig_125,sig_127,sig_136,sig_137,sig_138,sig_139,sig_140,sig_141,sig_142,sig_143,sig_144,sig_145;
wire sig_146,sig_147,sig_148,sig_149,sig_150,sig_151,sig_152,sig_153,sig_154,sig_155,sig_160,sig_162,sig_167,sig_169,sig_170,sig_171,sig_173,sig_175,sig_179,sig_184;
wire sig_186,sig_187,sig_189,sig_202,sig_204,sig_206,sig_208,sig_209,sig_210,sig_211,sig_212,sig_213,sig_215,sig_217,sig_221,sig_226,sig_227,sig_228,sig_229,sig_231;
wire sig_240,sig_241,sig_242,sig_243,sig_244,sig_245,sig_246,sig_247,sig_248,sig_249,sig_250,sig_251,sig_252,sig_253,sig_254,sig_255,sig_256,sig_257,sig_258,sig_259;
wire sig_264,sig_266,sig_271,sig_273,sig_274,sig_275,sig_277,sig_279,sig_283,sig_288,sig_290,sig_291,sig_293,sig_306,sig_308,sig_310,sig_312,sig_313,sig_314,sig_315;
wire sig_316,sig_317,sig_319,sig_321,sig_325,sig_330,sig_331,sig_332,sig_333,sig_335,sig_344,sig_345,sig_346,sig_347,sig_348,sig_349,sig_350,sig_351,sig_352,sig_353;
wire sig_354,sig_355,sig_356,sig_357,sig_358,sig_359,sig_360,sig_361,sig_362,sig_363,sig_368,sig_370,sig_375,sig_377,sig_378,sig_379,sig_381,sig_383,sig_387,sig_392;
wire sig_394,sig_395,sig_397,sig_410,sig_412,sig_414,sig_416,sig_417,sig_418,sig_419,sig_420,sig_421,sig_423,sig_425,sig_429,sig_434,sig_435,sig_436,sig_437,sig_439;
wire sig_460,sig_462,sig_464,sig_466,sig_467,sig_468,sig_469,sig_470,sig_471,sig_472,sig_473,sig_474,sig_475,sig_476,sig_477,sig_478,sig_479,sig_480,sig_481,sig_482;
wire sig_483,sig_484,sig_485,sig_486,sig_487,sig_488,sig_489,sig_490,sig_491,sig_492,sig_494,sig_499,sig_502,sig_506,sig_509,sig_510,sig_511,sig_512,sig_515,sig_516;
wire sig_517,sig_519,sig_520,sig_521,sig_550,sig_552,sig_554,sig_556,sig_557,sig_558,sig_559,sig_560,sig_561,sig_562,sig_563,sig_564,sig_565,sig_566,sig_567,sig_568;
wire sig_569,sig_570,sig_571,sig_572,sig_573,sig_574,sig_575,sig_576,sig_577,sig_578,sig_579,sig_580,sig_581,sig_582,sig_584,sig_589,sig_592,sig_596,sig_599,sig_600;
wire sig_601,sig_602,sig_605,sig_606,sig_607,sig_609,sig_610,sig_611,sig_628,sig_629,sig_630,sig_631,sig_632,sig_633,sig_634,sig_635,sig_636,sig_637,sig_638,sig_639;
wire sig_640,sig_641,sig_642,sig_643,sig_644,sig_645,sig_646,sig_647,sig_652,sig_654,sig_659,sig_661,sig_662,sig_663,sig_665,sig_667,sig_671,sig_676,sig_678,sig_679;
wire sig_681,sig_694,sig_696,sig_698,sig_700,sig_701,sig_702,sig_703,sig_704,sig_705,sig_707,sig_709,sig_713,sig_718,sig_719,sig_720,sig_721,sig_723,sig_732,sig_733;
wire sig_734,sig_735,sig_736,sig_737,sig_738,sig_739,sig_740,sig_741,sig_742,sig_743,sig_744,sig_745,sig_746,sig_747,sig_748,sig_749,sig_750,sig_751,sig_756,sig_758;
wire sig_763,sig_765,sig_766,sig_767,sig_769,sig_771,sig_775,sig_780,sig_782,sig_783,sig_785,sig_798,sig_800,sig_802,sig_804,sig_805,sig_806,sig_807,sig_808,sig_809;
wire sig_811,sig_813,sig_817,sig_822,sig_823,sig_824,sig_825,sig_827,sig_836,sig_837,sig_838,sig_839,sig_840,sig_841,sig_842,sig_843,sig_844,sig_845,sig_846,sig_847;
wire sig_848,sig_849,sig_850,sig_851,sig_852,sig_853,sig_854,sig_855,sig_860,sig_862,sig_867,sig_869,sig_870,sig_871,sig_873,sig_875,sig_879,sig_884,sig_886,sig_887;
wire sig_889,sig_902,sig_904,sig_906,sig_908,sig_909,sig_910,sig_911,sig_912,sig_913,sig_915,sig_917,sig_921,sig_926,sig_927,sig_928,sig_929,sig_931,sig_940,sig_941;
wire sig_942,sig_943,sig_944,sig_945,sig_946,sig_947,sig_948,sig_949,sig_950,sig_951,sig_952,sig_953,sig_954,sig_955,sig_956,sig_957,sig_958,sig_959,sig_964,sig_966;
wire sig_971,sig_973,sig_974,sig_975,sig_977,sig_979,sig_983,sig_988,sig_990,sig_991,sig_993,sig_1006,sig_1008,sig_1010,sig_1012,sig_1013,sig_1014,sig_1015,sig_1016,sig_1017;
wire sig_1019,sig_1021,sig_1025,sig_1030,sig_1031,sig_1032,sig_1033,sig_1035,sig_1056,sig_1058,sig_1060,sig_1062,sig_1063,sig_1064,sig_1065,sig_1066,sig_1067,sig_1068,sig_1069,sig_1070;
wire sig_1071,sig_1072,sig_1073,sig_1074,sig_1075,sig_1076,sig_1077,sig_1078,sig_1079,sig_1080,sig_1081,sig_1082,sig_1083,sig_1084,sig_1085,sig_1086,sig_1087,sig_1088,sig_1090,sig_1095;
wire sig_1098,sig_1102,sig_1105,sig_1106,sig_1107,sig_1108,sig_1111,sig_1112,sig_1113,sig_1115,sig_1116,sig_1117,sig_1146,sig_1148,sig_1150,sig_1152,sig_1153,sig_1154,sig_1155,sig_1156;
wire sig_1157,sig_1158,sig_1159,sig_1160,sig_1161,sig_1162,sig_1163,sig_1164,sig_1165,sig_1166,sig_1167,sig_1168,sig_1169,sig_1170,sig_1171,sig_1172,sig_1173,sig_1174,sig_1175,sig_1176;
wire sig_1177,sig_1178,sig_1180,sig_1185,sig_1188,sig_1192,sig_1195,sig_1196,sig_1197,sig_1198,sig_1201,sig_1202,sig_1203,sig_1205,sig_1206,sig_1207,sig_1224,sig_1225,sig_1226,sig_1227;
wire sig_1228,sig_1229,sig_1230,sig_1231,sig_1232,sig_1233,sig_1234,sig_1235,sig_1236,sig_1237,sig_1238,sig_1239,sig_1240,sig_1241,sig_1242,sig_1243,sig_1248,sig_1250,sig_1255,sig_1257;
wire sig_1258,sig_1259,sig_1261,sig_1263,sig_1267,sig_1272,sig_1274,sig_1275,sig_1277,sig_1290,sig_1292,sig_1294,sig_1296,sig_1297,sig_1298,sig_1299,sig_1300,sig_1301,sig_1303,sig_1305;
wire sig_1309,sig_1314,sig_1315,sig_1316,sig_1317,sig_1319,sig_1328,sig_1329,sig_1330,sig_1331,sig_1332,sig_1333,sig_1334,sig_1335,sig_1336,sig_1337,sig_1338,sig_1339,sig_1340,sig_1341;
wire sig_1342,sig_1343,sig_1344,sig_1345,sig_1346,sig_1347,sig_1352,sig_1354,sig_1359,sig_1361,sig_1362,sig_1363,sig_1365,sig_1367,sig_1371,sig_1376,sig_1378,sig_1379,sig_1381,sig_1394;
wire sig_1396,sig_1398,sig_1400,sig_1401,sig_1402,sig_1403,sig_1404,sig_1405,sig_1407,sig_1409,sig_1413,sig_1418,sig_1419,sig_1420,sig_1421,sig_1423,sig_1432,sig_1433,sig_1434,sig_1435;
wire sig_1436,sig_1437,sig_1438,sig_1439,sig_1440,sig_1441,sig_1442,sig_1443,sig_1444,sig_1445,sig_1446,sig_1447,sig_1448,sig_1449,sig_1450,sig_1451,sig_1456,sig_1458,sig_1463,sig_1465;
wire sig_1466,sig_1467,sig_1469,sig_1471,sig_1475,sig_1480,sig_1482,sig_1483,sig_1485,sig_1498,sig_1500,sig_1502,sig_1504,sig_1505,sig_1506,sig_1507,sig_1508,sig_1509,sig_1511,sig_1513;
wire sig_1517,sig_1522,sig_1523,sig_1524,sig_1525,sig_1527,sig_1536,sig_1537,sig_1538,sig_1539,sig_1540,sig_1541,sig_1542,sig_1543,sig_1544,sig_1545,sig_1546,sig_1547,sig_1548,sig_1549;
wire sig_1550,sig_1551,sig_1552,sig_1553,sig_1554,sig_1555,sig_1560,sig_1562,sig_1567,sig_1569,sig_1570,sig_1571,sig_1573,sig_1575,sig_1579,sig_1584,sig_1586,sig_1587,sig_1589,sig_1602;
wire sig_1604,sig_1606,sig_1608,sig_1609,sig_1610,sig_1611,sig_1612,sig_1613,sig_1615,sig_1617,sig_1621,sig_1626,sig_1627,sig_1628,sig_1629,sig_1631,sig_1652,sig_1654,sig_1656,sig_1658;
wire sig_1659,sig_1660,sig_1661,sig_1662,sig_1663,sig_1664,sig_1665,sig_1666,sig_1667,sig_1668,sig_1669,sig_1670,sig_1671,sig_1672,sig_1673,sig_1674,sig_1675,sig_1676,sig_1677,sig_1678;
wire sig_1679,sig_1680,sig_1681,sig_1682,sig_1683,sig_1684,sig_1686,sig_1691,sig_1694,sig_1698,sig_1701,sig_1702,sig_1703,sig_1704,sig_1707,sig_1708,sig_1709,sig_1711,sig_1712,sig_1713;
wire sig_1742,sig_1744,sig_1746,sig_1748,sig_1749,sig_1750,sig_1751,sig_1752,sig_1753,sig_1754,sig_1755,sig_1756,sig_1757,sig_1758,sig_1759,sig_1760,sig_1761,sig_1762,sig_1763,sig_1764;
wire sig_1765,sig_1766,sig_1767,sig_1768,sig_1769,sig_1770,sig_1771,sig_1772,sig_1773,sig_1774,sig_1776,sig_1781,sig_1784,sig_1788,sig_1791,sig_1792,sig_1793,sig_1794,sig_1797,sig_1798;
wire sig_1799,sig_1801,sig_1802,sig_1803,sig_1820,sig_1821,sig_1822,sig_1823,sig_1824,sig_1825,sig_1826,sig_1827,sig_1828,sig_1829,sig_1830,sig_1831,sig_1832,sig_1833,sig_1834,sig_1835;
wire sig_1836,sig_1837,sig_1838,sig_1839,sig_1844,sig_1846,sig_1851,sig_1853,sig_1854,sig_1855,sig_1857,sig_1859,sig_1863,sig_1868,sig_1870,sig_1871,sig_1873,sig_1886,sig_1888,sig_1890;
wire sig_1892,sig_1893,sig_1894,sig_1895,sig_1896,sig_1897,sig_1899,sig_1901,sig_1905,sig_1910,sig_1911,sig_1912,sig_1913,sig_1915,sig_1924,sig_1925,sig_1926,sig_1927,sig_1928,sig_1929;
wire sig_1930,sig_1931,sig_1932,sig_1933,sig_1934,sig_1935,sig_1936,sig_1937,sig_1938,sig_1939,sig_1940,sig_1941,sig_1942,sig_1943,sig_1948,sig_1950,sig_1955,sig_1957,sig_1958,sig_1959;
wire sig_1961,sig_1963,sig_1967,sig_1972,sig_1974,sig_1975,sig_1977,sig_1990,sig_1992,sig_1994,sig_1996,sig_1997,sig_1998,sig_1999,sig_2000,sig_2001,sig_2003,sig_2005,sig_2009,sig_2014;
wire sig_2015,sig_2016,sig_2017,sig_2019,sig_2028,sig_2029,sig_2030,sig_2031,sig_2032,sig_2033,sig_2034,sig_2035,sig_2036,sig_2037,sig_2038,sig_2039,sig_2040,sig_2041,sig_2042,sig_2043;
wire sig_2044,sig_2045,sig_2046,sig_2047,sig_2052,sig_2054,sig_2059,sig_2061,sig_2062,sig_2063,sig_2065,sig_2067,sig_2071,sig_2076,sig_2078,sig_2079,sig_2081,sig_2094,sig_2096,sig_2098;
wire sig_2100,sig_2101,sig_2102,sig_2103,sig_2104,sig_2105,sig_2107,sig_2109,sig_2113,sig_2118,sig_2119,sig_2120,sig_2121,sig_2123,sig_2132,sig_2133,sig_2134,sig_2135,sig_2136,sig_2137;
wire sig_2138,sig_2139,sig_2140,sig_2141,sig_2142,sig_2143,sig_2144,sig_2145,sig_2146,sig_2147,sig_2148,sig_2149,sig_2150,sig_2151,sig_2156,sig_2158,sig_2163,sig_2165,sig_2166,sig_2167;
wire sig_2169,sig_2171,sig_2175,sig_2180,sig_2182,sig_2183,sig_2185,sig_2198,sig_2200,sig_2202,sig_2204,sig_2205,sig_2206,sig_2207,sig_2208,sig_2209,sig_2211,sig_2213,sig_2217,sig_2222;
wire sig_2223,sig_2224,sig_2225,sig_2227,sig_2248,sig_2250,sig_2252,sig_2254,sig_2255,sig_2256,sig_2257,sig_2258,sig_2259,sig_2260,sig_2261,sig_2262,sig_2263,sig_2264,sig_2265,sig_2266;
wire sig_2267,sig_2268,sig_2269,sig_2270,sig_2271,sig_2272,sig_2273,sig_2274,sig_2275,sig_2276,sig_2277,sig_2278,sig_2279,sig_2280,sig_2282,sig_2287,sig_2290,sig_2294,sig_2297,sig_2298;
wire sig_2299,sig_2300,sig_2303,sig_2304,sig_2305,sig_2307,sig_2308,sig_2309,sig_2338,sig_2340,sig_2342,sig_2344,sig_2345,sig_2346,sig_2347,sig_2348,sig_2349,sig_2350,sig_2351,sig_2352;
wire sig_2353,sig_2354,sig_2355,sig_2356,sig_2357,sig_2358,sig_2359,sig_2360,sig_2361,sig_2362,sig_2363,sig_2364,sig_2365,sig_2366,sig_2367,sig_2368,sig_2369,sig_2370,sig_2372,sig_2377;
wire sig_2380,sig_2384,sig_2387,sig_2388,sig_2389,sig_2390,sig_2393,sig_2394,sig_2395,sig_2397,sig_2398,sig_2399,sig_2432,sig_2433,sig_2434,sig_2435,sig_2436,sig_2437,sig_2438,sig_2439;
wire sig_2440,sig_2441,sig_2442,sig_2443,sig_2444,sig_2445,sig_2446,sig_2447,sig_2448,sig_2449,sig_2450,sig_2451,sig_2452,sig_2453,sig_2454,sig_2455,sig_2456,sig_2457,sig_2458,sig_2459;
wire sig_2460,sig_2461,sig_2462,sig_2463,sig_2503,sig_2504,sig_2505,sig_2506,sig_2507,sig_2508,sig_2509,sig_2510,sig_2511,sig_2512,sig_2513,sig_2514,sig_2515,sig_2516,sig_2517,sig_2518;
wire sig_2519,sig_2520,sig_2521,sig_2522,sig_2523,sig_2524,sig_2525,sig_2526,sig_2527,sig_2528,sig_2529,sig_2530,sig_2531,sig_2532,sig_2533,sig_2534,sig_2535,sig_2536,sig_2537,sig_2538;
wire sig_2539,sig_2540,sig_2541,sig_2542,sig_2543,sig_2544,sig_2545,sig_2546,sig_2547,sig_2548,sig_2549,sig_2551,sig_2552,sig_2554,sig_2555,sig_2557,sig_2558,sig_2560,sig_2561,sig_2563;
wire sig_2564,sig_2566,sig_2567,sig_2569,sig_2586,sig_2587,sig_2588,sig_2589,sig_2590,sig_2591,sig_2592,sig_2593,sig_2594,sig_2595,sig_2596,sig_2597,sig_2598,sig_2599,sig_2600,sig_2601;
wire sig_2602,sig_2603,sig_2604,sig_2605,sig_2606,sig_2607,sig_2608,sig_2609,sig_2610,sig_2611,sig_2612,sig_2613,sig_2614,sig_2615,sig_2616,sig_2617,sig_2657,sig_2658,sig_2659,sig_2660;
wire sig_2661,sig_2662,sig_2663,sig_2664,sig_2665,sig_2666,sig_2667,sig_2668,sig_2669,sig_2670,sig_2671,sig_2672,sig_2673,sig_2674,sig_2675,sig_2676,sig_2677,sig_2678,sig_2679,sig_2680;
wire sig_2681,sig_2682,sig_2683,sig_2684,sig_2685,sig_2686,sig_2687,sig_2688,sig_2689,sig_2690,sig_2691,sig_2692,sig_2693,sig_2694,sig_2695,sig_2696,sig_2697,sig_2698,sig_2699,sig_2700;
wire sig_2701,sig_2702,sig_2703,sig_2705,sig_2706,sig_2708,sig_2709,sig_2711,sig_2712,sig_2714,sig_2715,sig_2717,sig_2718,sig_2720,sig_2721,sig_2723;

assign sig_32 = A[1] & B[0];
assign sig_33 = A[1] & B[1];
assign sig_34 = B[1] & A[0];
assign sig_35 = A[0] & B[0];
assign sig_36 = sig_34 | sig_32;
assign sig_37 = A[3] & B[0];
assign sig_38 = A[3] & B[1];
assign sig_39 = B[1] & A[2];
assign sig_40 = A[2] & B[0];
assign sig_41 = sig_39 | sig_37;
assign sig_42 = A[1] & B[2];
assign sig_43 = A[1] & B[3];
assign sig_44 = B[3] & A[0];
assign sig_45 = A[0] & B[2];
assign sig_46 = sig_44 | sig_42;
assign sig_47 = A[3] & B[2];
assign sig_48 = A[3] & B[3];
assign sig_49 = B[3] & A[2];
assign sig_50 = A[2] & B[2];
assign sig_51 = sig_49 | sig_47;
assign sig_56 = sig_40 ^ sig_33;
assign sig_58 = sig_40 & sig_33;
assign sig_63 = sig_41 & sig_58;
assign sig_65 = sig_38 ^ sig_50;
assign sig_66 = sig_38 & sig_50;
assign sig_67 = sig_65 & sig_63;
assign sig_69 = sig_66 | sig_67;
assign sig_71 = sig_51 & sig_69;
assign sig_75 = sig_48 & sig_71;
assign sig_80 = sig_65 ^ sig_63;
assign sig_82 = sig_48 ^ sig_71;
assign sig_83 = sig_51 ^ sig_69;
assign sig_85 = sig_41 ^ sig_58;
assign sig_98 = sig_45 ^ sig_56;
assign sig_100 = sig_45 & sig_56;
assign sig_102 = sig_46 ^ sig_85;
assign sig_104 = sig_46 & sig_85;
assign sig_105 = sig_102 & sig_100;
assign sig_106 = sig_104 | sig_105;
assign sig_107 = sig_43 ^ sig_80;
assign sig_108 = sig_43 & sig_80;
assign sig_109 = sig_107 & sig_106;
assign sig_111 = sig_108 | sig_109;
assign sig_113 = sig_83 & sig_111;
assign sig_117 = sig_82 & sig_113;
assign sig_122 = sig_107 ^ sig_106;
assign sig_123 = sig_75 ^ sig_117;
assign sig_124 = sig_82 ^ sig_113;
assign sig_125 = sig_83 ^ sig_111;
assign sig_127 = sig_102 ^ sig_100;
assign sig_136 = A[5] & B[0];
assign sig_137 = A[5] & B[1];
assign sig_138 = B[1] & A[4];
assign sig_139 = A[4] & B[0];
assign sig_140 = sig_138 | sig_136;
assign sig_141 = A[7] & B[0];
assign sig_142 = A[7] & B[1];
assign sig_143 = B[1] & A[6];
assign sig_144 = A[6] & B[0];
assign sig_145 = sig_143 | sig_141;
assign sig_146 = A[5] & B[2];
assign sig_147 = A[5] & B[3];
assign sig_148 = B[3] & A[4];
assign sig_149 = A[4] & B[2];
assign sig_150 = sig_148 | sig_146;
assign sig_151 = A[7] & B[2];
assign sig_152 = A[7] & B[3];
assign sig_153 = B[3] & A[6];
assign sig_154 = A[6] & B[2];
assign sig_155 = sig_153 | sig_151;
assign sig_160 = sig_144 ^ sig_137;
assign sig_162 = sig_144 & sig_137;
assign sig_167 = sig_145 & sig_162;
assign sig_169 = sig_142 ^ sig_154;
assign sig_170 = sig_142 & sig_154;
assign sig_171 = sig_169 & sig_167;
assign sig_173 = sig_170 | sig_171;
assign sig_175 = sig_155 & sig_173;
assign sig_179 = sig_152 & sig_175;
assign sig_184 = sig_169 ^ sig_167;
assign sig_186 = sig_152 ^ sig_175;
assign sig_187 = sig_155 ^ sig_173;
assign sig_189 = sig_145 ^ sig_162;
assign sig_202 = sig_149 ^ sig_160;
assign sig_204 = sig_149 & sig_160;
assign sig_206 = sig_150 ^ sig_189;
assign sig_208 = sig_150 & sig_189;
assign sig_209 = sig_206 & sig_204;
assign sig_210 = sig_208 | sig_209;
assign sig_211 = sig_147 ^ sig_184;
assign sig_212 = sig_147 & sig_184;
assign sig_213 = sig_211 & sig_210;
assign sig_215 = sig_212 | sig_213;
assign sig_217 = sig_187 & sig_215;
assign sig_221 = sig_186 & sig_217;
assign sig_226 = sig_211 ^ sig_210;
assign sig_227 = sig_179 ^ sig_221;
assign sig_228 = sig_186 ^ sig_217;
assign sig_229 = sig_187 ^ sig_215;
assign sig_231 = sig_206 ^ sig_204;
assign sig_240 = A[1] & B[4];
assign sig_241 = A[1] & B[5];
assign sig_242 = B[5] & A[0];
assign sig_243 = A[0] & B[4];
assign sig_244 = sig_242 | sig_240;
assign sig_245 = A[3] & B[4];
assign sig_246 = A[3] & B[5];
assign sig_247 = B[5] & A[2];
assign sig_248 = A[2] & B[4];
assign sig_249 = sig_247 | sig_245;
assign sig_250 = A[1] & B[6];
assign sig_251 = A[1] & B[7];
assign sig_252 = B[7] & A[0];
assign sig_253 = A[0] & B[6];
assign sig_254 = sig_252 | sig_250;
assign sig_255 = A[3] & B[6];
assign sig_256 = A[3] & B[7];
assign sig_257 = B[7] & A[2];
assign sig_258 = A[2] & B[6];
assign sig_259 = sig_257 | sig_255;
assign sig_264 = sig_248 ^ sig_241;
assign sig_266 = sig_248 & sig_241;
assign sig_271 = sig_249 & sig_266;
assign sig_273 = sig_246 ^ sig_258;
assign sig_274 = sig_246 & sig_258;
assign sig_275 = sig_273 & sig_271;
assign sig_277 = sig_274 | sig_275;
assign sig_279 = sig_259 & sig_277;
assign sig_283 = sig_256 & sig_279;
assign sig_288 = sig_273 ^ sig_271;
assign sig_290 = sig_256 ^ sig_279;
assign sig_291 = sig_259 ^ sig_277;
assign sig_293 = sig_249 ^ sig_266;
assign sig_306 = sig_253 ^ sig_264;
assign sig_308 = sig_253 & sig_264;
assign sig_310 = sig_254 ^ sig_293;
assign sig_312 = sig_254 & sig_293;
assign sig_313 = sig_310 & sig_308;
assign sig_314 = sig_312 | sig_313;
assign sig_315 = sig_251 ^ sig_288;
assign sig_316 = sig_251 & sig_288;
assign sig_317 = sig_315 & sig_314;
assign sig_319 = sig_316 | sig_317;
assign sig_321 = sig_291 & sig_319;
assign sig_325 = sig_290 & sig_321;
assign sig_330 = sig_315 ^ sig_314;
assign sig_331 = sig_283 ^ sig_325;
assign sig_332 = sig_290 ^ sig_321;
assign sig_333 = sig_291 ^ sig_319;
assign sig_335 = sig_310 ^ sig_308;
assign sig_344 = A[5] & B[4];
assign sig_345 = A[5] & B[5];
assign sig_346 = B[5] & A[4];
assign sig_347 = A[4] & B[4];
assign sig_348 = sig_346 | sig_344;
assign sig_349 = A[7] & B[4];
assign sig_350 = A[7] & B[5];
assign sig_351 = B[5] & A[6];
assign sig_352 = A[6] & B[4];
assign sig_353 = sig_351 | sig_349;
assign sig_354 = A[5] & B[6];
assign sig_355 = A[5] & B[7];
assign sig_356 = B[7] & A[4];
assign sig_357 = A[4] & B[6];
assign sig_358 = sig_356 | sig_354;
assign sig_359 = A[7] & B[6];
assign sig_360 = A[7] & B[7];
assign sig_361 = B[7] & A[6];
assign sig_362 = A[6] & B[6];
assign sig_363 = sig_361 | sig_359;
assign sig_368 = sig_352 ^ sig_345;
assign sig_370 = sig_352 & sig_345;
assign sig_375 = sig_353 & sig_370;
assign sig_377 = sig_350 ^ sig_362;
assign sig_378 = sig_350 & sig_362;
assign sig_379 = sig_377 & sig_375;
assign sig_381 = sig_378 | sig_379;
assign sig_383 = sig_363 & sig_381;
assign sig_387 = sig_360 & sig_383;
assign sig_392 = sig_377 ^ sig_375;
assign sig_394 = sig_360 ^ sig_383;
assign sig_395 = sig_363 ^ sig_381;
assign sig_397 = sig_353 ^ sig_370;
assign sig_410 = sig_357 ^ sig_368;
assign sig_412 = sig_357 & sig_368;
assign sig_414 = sig_358 ^ sig_397;
assign sig_416 = sig_358 & sig_397;
assign sig_417 = sig_414 & sig_412;
assign sig_418 = sig_416 | sig_417;
assign sig_419 = sig_355 ^ sig_392;
assign sig_420 = sig_355 & sig_392;
assign sig_421 = sig_419 & sig_418;
assign sig_423 = sig_420 | sig_421;
assign sig_425 = sig_395 & sig_423;
assign sig_429 = sig_394 & sig_425;
assign sig_434 = sig_419 ^ sig_418;
assign sig_435 = sig_387 ^ sig_429;
assign sig_436 = sig_394 ^ sig_425;
assign sig_437 = sig_395 ^ sig_423;
assign sig_439 = sig_414 ^ sig_412;
assign sig_460 = sig_139 ^ sig_122;
assign sig_462 = sig_139 & sig_122;
assign sig_464 = sig_140 ^ sig_125;
assign sig_466 = sig_464 & sig_462;
assign sig_467 = sig_140 & sig_125;
assign sig_468 = sig_467 | sig_466;
assign sig_469 = sig_202 ^ sig_124;
assign sig_470 = sig_469 & sig_468;
assign sig_471 = sig_202 & sig_124;
assign sig_472 = sig_471 | sig_470;
assign sig_473 = sig_231 ^ sig_123;
assign sig_474 = sig_473 & sig_472;
assign sig_475 = sig_231 & sig_123;
assign sig_476 = sig_226 ^ sig_347;
assign sig_477 = sig_475 | sig_474;
assign sig_478 = sig_226 & sig_347;
assign sig_479 = sig_476 & sig_477;
assign sig_480 = sig_229 ^ sig_348;
assign sig_481 = sig_478 | sig_479;
assign sig_482 = sig_229 & sig_348;
assign sig_483 = sig_480 & sig_481;
assign sig_484 = sig_228 ^ sig_410;
assign sig_485 = sig_482 | sig_483;
assign sig_486 = sig_484 & sig_485;
assign sig_487 = sig_228 & sig_410;
assign sig_488 = sig_487 | sig_486;
assign sig_489 = sig_227 ^ sig_439;
assign sig_490 = sig_489 & sig_488;
assign sig_491 = sig_227 & sig_439;
assign sig_492 = sig_491 | sig_490;
assign sig_494 = sig_434 & sig_492;
assign sig_499 = sig_437 & sig_494;
assign sig_502 = sig_436 & sig_499;
assign sig_506 = sig_464 ^ sig_462;
assign sig_509 = sig_484 ^ sig_485;
assign sig_510 = sig_469 ^ sig_468;
assign sig_511 = sig_489 ^ sig_488;
assign sig_512 = sig_434 ^ sig_492;
assign sig_515 = sig_437 ^ sig_494;
assign sig_516 = sig_436 ^ sig_499;
assign sig_517 = sig_480 ^ sig_481;
assign sig_519 = sig_435 ^ sig_502;
assign sig_520 = sig_476 ^ sig_477;
assign sig_521 = sig_473 ^ sig_472;
assign sig_550 = sig_243 ^ sig_460;
assign sig_552 = sig_243 & sig_460;
assign sig_554 = sig_244 ^ sig_506;
assign sig_556 = sig_554 & sig_552;
assign sig_557 = sig_244 & sig_506;
assign sig_558 = sig_557 | sig_556;
assign sig_559 = sig_306 ^ sig_510;
assign sig_560 = sig_559 & sig_558;
assign sig_561 = sig_306 & sig_510;
assign sig_562 = sig_561 | sig_560;
assign sig_563 = sig_335 ^ sig_521;
assign sig_564 = sig_563 & sig_562;
assign sig_565 = sig_335 & sig_521;
assign sig_566 = sig_330 ^ sig_520;
assign sig_567 = sig_565 | sig_564;
assign sig_568 = sig_330 & sig_520;
assign sig_569 = sig_566 & sig_567;
assign sig_570 = sig_333 ^ sig_517;
assign sig_571 = sig_568 | sig_569;
assign sig_572 = sig_333 & sig_517;
assign sig_573 = sig_570 & sig_571;
assign sig_574 = sig_332 ^ sig_509;
assign sig_575 = sig_572 | sig_573;
assign sig_576 = sig_574 & sig_575;
assign sig_577 = sig_332 & sig_509;
assign sig_578 = sig_577 | sig_576;
assign sig_579 = sig_331 ^ sig_511;
assign sig_580 = sig_579 & sig_578;
assign sig_581 = sig_331 & sig_511;
assign sig_582 = sig_581 | sig_580;
assign sig_584 = sig_512 & sig_582;
assign sig_589 = sig_515 & sig_584;
assign sig_592 = sig_516 & sig_589;
assign sig_596 = sig_554 ^ sig_552;
assign sig_599 = sig_574 ^ sig_575;
assign sig_600 = sig_559 ^ sig_558;
assign sig_601 = sig_579 ^ sig_578;
assign sig_602 = sig_512 ^ sig_582;
assign sig_605 = sig_515 ^ sig_584;
assign sig_606 = sig_516 ^ sig_589;
assign sig_607 = sig_570 ^ sig_571;
assign sig_609 = sig_519 ^ sig_592;
assign sig_610 = sig_566 ^ sig_567;
assign sig_611 = sig_563 ^ sig_562;
assign sig_628 = A[9] & B[0];
assign sig_629 = A[9] & B[1];
assign sig_630 = B[1] & A[8];
assign sig_631 = A[8] & B[0];
assign sig_632 = sig_630 | sig_628;
assign sig_633 = A[11] & B[0];
assign sig_634 = A[11] & B[1];
assign sig_635 = B[1] & A[10];
assign sig_636 = A[10] & B[0];
assign sig_637 = sig_635 | sig_633;
assign sig_638 = A[9] & B[2];
assign sig_639 = A[9] & B[3];
assign sig_640 = B[3] & A[8];
assign sig_641 = A[8] & B[2];
assign sig_642 = sig_640 | sig_638;
assign sig_643 = A[11] & B[2];
assign sig_644 = A[11] & B[3];
assign sig_645 = B[3] & A[10];
assign sig_646 = A[10] & B[2];
assign sig_647 = sig_645 | sig_643;
assign sig_652 = sig_636 ^ sig_629;
assign sig_654 = sig_636 & sig_629;
assign sig_659 = sig_637 & sig_654;
assign sig_661 = sig_634 ^ sig_646;
assign sig_662 = sig_634 & sig_646;
assign sig_663 = sig_661 & sig_659;
assign sig_665 = sig_662 | sig_663;
assign sig_667 = sig_647 & sig_665;
assign sig_671 = sig_644 & sig_667;
assign sig_676 = sig_661 ^ sig_659;
assign sig_678 = sig_644 ^ sig_667;
assign sig_679 = sig_647 ^ sig_665;
assign sig_681 = sig_637 ^ sig_654;
assign sig_694 = sig_641 ^ sig_652;
assign sig_696 = sig_641 & sig_652;
assign sig_698 = sig_642 ^ sig_681;
assign sig_700 = sig_642 & sig_681;
assign sig_701 = sig_698 & sig_696;
assign sig_702 = sig_700 | sig_701;
assign sig_703 = sig_639 ^ sig_676;
assign sig_704 = sig_639 & sig_676;
assign sig_705 = sig_703 & sig_702;
assign sig_707 = sig_704 | sig_705;
assign sig_709 = sig_679 & sig_707;
assign sig_713 = sig_678 & sig_709;
assign sig_718 = sig_703 ^ sig_702;
assign sig_719 = sig_671 ^ sig_713;
assign sig_720 = sig_678 ^ sig_709;
assign sig_721 = sig_679 ^ sig_707;
assign sig_723 = sig_698 ^ sig_696;
assign sig_732 = A[13] & B[0];
assign sig_733 = A[13] & B[1];
assign sig_734 = B[1] & A[12];
assign sig_735 = A[12] & B[0];
assign sig_736 = sig_734 | sig_732;
assign sig_737 = A[15] & B[0];
assign sig_738 = A[15] & B[1];
assign sig_739 = B[1] & A[14];
assign sig_740 = A[14] & B[0];
assign sig_741 = sig_739 | sig_737;
assign sig_742 = A[13] & B[2];
assign sig_743 = A[13] & B[3];
assign sig_744 = B[3] & A[12];
assign sig_745 = A[12] & B[2];
assign sig_746 = sig_744 | sig_742;
assign sig_747 = A[15] & B[2];
assign sig_748 = A[15] & B[3];
assign sig_749 = B[3] & A[14];
assign sig_750 = A[14] & B[2];
assign sig_751 = sig_749 | sig_747;
assign sig_756 = sig_740 ^ sig_733;
assign sig_758 = sig_740 & sig_733;
assign sig_763 = sig_741 & sig_758;
assign sig_765 = sig_738 ^ sig_750;
assign sig_766 = sig_738 & sig_750;
assign sig_767 = sig_765 & sig_763;
assign sig_769 = sig_766 | sig_767;
assign sig_771 = sig_751 & sig_769;
assign sig_775 = sig_748 & sig_771;
assign sig_780 = sig_765 ^ sig_763;
assign sig_782 = sig_748 ^ sig_771;
assign sig_783 = sig_751 ^ sig_769;
assign sig_785 = sig_741 ^ sig_758;
assign sig_798 = sig_745 ^ sig_756;
assign sig_800 = sig_745 & sig_756;
assign sig_802 = sig_746 ^ sig_785;
assign sig_804 = sig_746 & sig_785;
assign sig_805 = sig_802 & sig_800;
assign sig_806 = sig_804 | sig_805;
assign sig_807 = sig_743 ^ sig_780;
assign sig_808 = sig_743 & sig_780;
assign sig_809 = sig_807 & sig_806;
assign sig_811 = sig_808 | sig_809;
assign sig_813 = sig_783 & sig_811;
assign sig_817 = sig_782 & sig_813;
assign sig_822 = sig_807 ^ sig_806;
assign sig_823 = sig_775 ^ sig_817;
assign sig_824 = sig_782 ^ sig_813;
assign sig_825 = sig_783 ^ sig_811;
assign sig_827 = sig_802 ^ sig_800;
assign sig_836 = A[9] & B[4];
assign sig_837 = A[9] & B[5];
assign sig_838 = B[5] & A[8];
assign sig_839 = A[8] & B[4];
assign sig_840 = sig_838 | sig_836;
assign sig_841 = A[11] & B[4];
assign sig_842 = A[11] & B[5];
assign sig_843 = B[5] & A[10];
assign sig_844 = A[10] & B[4];
assign sig_845 = sig_843 | sig_841;
assign sig_846 = A[9] & B[6];
assign sig_847 = A[9] & B[7];
assign sig_848 = B[7] & A[8];
assign sig_849 = A[8] & B[6];
assign sig_850 = sig_848 | sig_846;
assign sig_851 = A[11] & B[6];
assign sig_852 = A[11] & B[7];
assign sig_853 = B[7] & A[10];
assign sig_854 = A[10] & B[6];
assign sig_855 = sig_853 | sig_851;
assign sig_860 = sig_844 ^ sig_837;
assign sig_862 = sig_844 & sig_837;
assign sig_867 = sig_845 & sig_862;
assign sig_869 = sig_842 ^ sig_854;
assign sig_870 = sig_842 & sig_854;
assign sig_871 = sig_869 & sig_867;
assign sig_873 = sig_870 | sig_871;
assign sig_875 = sig_855 & sig_873;
assign sig_879 = sig_852 & sig_875;
assign sig_884 = sig_869 ^ sig_867;
assign sig_886 = sig_852 ^ sig_875;
assign sig_887 = sig_855 ^ sig_873;
assign sig_889 = sig_845 ^ sig_862;
assign sig_902 = sig_849 ^ sig_860;
assign sig_904 = sig_849 & sig_860;
assign sig_906 = sig_850 ^ sig_889;
assign sig_908 = sig_850 & sig_889;
assign sig_909 = sig_906 & sig_904;
assign sig_910 = sig_908 | sig_909;
assign sig_911 = sig_847 ^ sig_884;
assign sig_912 = sig_847 & sig_884;
assign sig_913 = sig_911 & sig_910;
assign sig_915 = sig_912 | sig_913;
assign sig_917 = sig_887 & sig_915;
assign sig_921 = sig_886 & sig_917;
assign sig_926 = sig_911 ^ sig_910;
assign sig_927 = sig_879 ^ sig_921;
assign sig_928 = sig_886 ^ sig_917;
assign sig_929 = sig_887 ^ sig_915;
assign sig_931 = sig_906 ^ sig_904;
assign sig_940 = A[13] & B[4];
assign sig_941 = A[13] & B[5];
assign sig_942 = B[5] & A[12];
assign sig_943 = A[12] & B[4];
assign sig_944 = sig_942 | sig_940;
assign sig_945 = A[15] & B[4];
assign sig_946 = A[15] & B[5];
assign sig_947 = B[5] & A[14];
assign sig_948 = A[14] & B[4];
assign sig_949 = sig_947 | sig_945;
assign sig_950 = A[13] & B[6];
assign sig_951 = A[13] & B[7];
assign sig_952 = B[7] & A[12];
assign sig_953 = A[12] & B[6];
assign sig_954 = sig_952 | sig_950;
assign sig_955 = A[15] & B[6];
assign sig_956 = A[15] & B[7];
assign sig_957 = B[7] & A[14];
assign sig_958 = A[14] & B[6];
assign sig_959 = sig_957 | sig_955;
assign sig_964 = sig_948 ^ sig_941;
assign sig_966 = sig_948 & sig_941;
assign sig_971 = sig_949 & sig_966;
assign sig_973 = sig_946 ^ sig_958;
assign sig_974 = sig_946 & sig_958;
assign sig_975 = sig_973 & sig_971;
assign sig_977 = sig_974 | sig_975;
assign sig_979 = sig_959 & sig_977;
assign sig_983 = sig_956 & sig_979;
assign sig_988 = sig_973 ^ sig_971;
assign sig_990 = sig_956 ^ sig_979;
assign sig_991 = sig_959 ^ sig_977;
assign sig_993 = sig_949 ^ sig_966;
assign sig_1006 = sig_953 ^ sig_964;
assign sig_1008 = sig_953 & sig_964;
assign sig_1010 = sig_954 ^ sig_993;
assign sig_1012 = sig_954 & sig_993;
assign sig_1013 = sig_1010 & sig_1008;
assign sig_1014 = sig_1012 | sig_1013;
assign sig_1015 = sig_951 ^ sig_988;
assign sig_1016 = sig_951 & sig_988;
assign sig_1017 = sig_1015 & sig_1014;
assign sig_1019 = sig_1016 | sig_1017;
assign sig_1021 = sig_991 & sig_1019;
assign sig_1025 = sig_990 & sig_1021;
assign sig_1030 = sig_1015 ^ sig_1014;
assign sig_1031 = sig_983 ^ sig_1025;
assign sig_1032 = sig_990 ^ sig_1021;
assign sig_1033 = sig_991 ^ sig_1019;
assign sig_1035 = sig_1010 ^ sig_1008;
assign sig_1056 = sig_735 ^ sig_718;
assign sig_1058 = sig_735 & sig_718;
assign sig_1060 = sig_736 ^ sig_721;
assign sig_1062 = sig_1060 & sig_1058;
assign sig_1063 = sig_736 & sig_721;
assign sig_1064 = sig_1063 | sig_1062;
assign sig_1065 = sig_798 ^ sig_720;
assign sig_1066 = sig_1065 & sig_1064;
assign sig_1067 = sig_798 & sig_720;
assign sig_1068 = sig_1067 | sig_1066;
assign sig_1069 = sig_827 ^ sig_719;
assign sig_1070 = sig_1069 & sig_1068;
assign sig_1071 = sig_827 & sig_719;
assign sig_1072 = sig_822 ^ sig_943;
assign sig_1073 = sig_1071 | sig_1070;
assign sig_1074 = sig_822 & sig_943;
assign sig_1075 = sig_1072 & sig_1073;
assign sig_1076 = sig_825 ^ sig_944;
assign sig_1077 = sig_1074 | sig_1075;
assign sig_1078 = sig_825 & sig_944;
assign sig_1079 = sig_1076 & sig_1077;
assign sig_1080 = sig_824 ^ sig_1006;
assign sig_1081 = sig_1078 | sig_1079;
assign sig_1082 = sig_1080 & sig_1081;
assign sig_1083 = sig_824 & sig_1006;
assign sig_1084 = sig_1083 | sig_1082;
assign sig_1085 = sig_823 ^ sig_1035;
assign sig_1086 = sig_1085 & sig_1084;
assign sig_1087 = sig_823 & sig_1035;
assign sig_1088 = sig_1087 | sig_1086;
assign sig_1090 = sig_1030 & sig_1088;
assign sig_1095 = sig_1033 & sig_1090;
assign sig_1098 = sig_1032 & sig_1095;
assign sig_1102 = sig_1060 ^ sig_1058;
assign sig_1105 = sig_1080 ^ sig_1081;
assign sig_1106 = sig_1065 ^ sig_1064;
assign sig_1107 = sig_1085 ^ sig_1084;
assign sig_1108 = sig_1030 ^ sig_1088;
assign sig_1111 = sig_1033 ^ sig_1090;
assign sig_1112 = sig_1032 ^ sig_1095;
assign sig_1113 = sig_1076 ^ sig_1077;
assign sig_1115 = sig_1031 ^ sig_1098;
assign sig_1116 = sig_1072 ^ sig_1073;
assign sig_1117 = sig_1069 ^ sig_1068;
assign sig_1146 = sig_839 ^ sig_1056;
assign sig_1148 = sig_839 & sig_1056;
assign sig_1150 = sig_840 ^ sig_1102;
assign sig_1152 = sig_1150 & sig_1148;
assign sig_1153 = sig_840 & sig_1102;
assign sig_1154 = sig_1153 | sig_1152;
assign sig_1155 = sig_902 ^ sig_1106;
assign sig_1156 = sig_1155 & sig_1154;
assign sig_1157 = sig_902 & sig_1106;
assign sig_1158 = sig_1157 | sig_1156;
assign sig_1159 = sig_931 ^ sig_1117;
assign sig_1160 = sig_1159 & sig_1158;
assign sig_1161 = sig_931 & sig_1117;
assign sig_1162 = sig_926 ^ sig_1116;
assign sig_1163 = sig_1161 | sig_1160;
assign sig_1164 = sig_926 & sig_1116;
assign sig_1165 = sig_1162 & sig_1163;
assign sig_1166 = sig_929 ^ sig_1113;
assign sig_1167 = sig_1164 | sig_1165;
assign sig_1168 = sig_929 & sig_1113;
assign sig_1169 = sig_1166 & sig_1167;
assign sig_1170 = sig_928 ^ sig_1105;
assign sig_1171 = sig_1168 | sig_1169;
assign sig_1172 = sig_1170 & sig_1171;
assign sig_1173 = sig_928 & sig_1105;
assign sig_1174 = sig_1173 | sig_1172;
assign sig_1175 = sig_927 ^ sig_1107;
assign sig_1176 = sig_1175 & sig_1174;
assign sig_1177 = sig_927 & sig_1107;
assign sig_1178 = sig_1177 | sig_1176;
assign sig_1180 = sig_1108 & sig_1178;
assign sig_1185 = sig_1111 & sig_1180;
assign sig_1188 = sig_1112 & sig_1185;
assign sig_1192 = sig_1150 ^ sig_1148;
assign sig_1195 = sig_1170 ^ sig_1171;
assign sig_1196 = sig_1155 ^ sig_1154;
assign sig_1197 = sig_1175 ^ sig_1174;
assign sig_1198 = sig_1108 ^ sig_1178;
assign sig_1201 = sig_1111 ^ sig_1180;
assign sig_1202 = sig_1112 ^ sig_1185;
assign sig_1203 = sig_1166 ^ sig_1167;
assign sig_1205 = sig_1115 ^ sig_1188;
assign sig_1206 = sig_1162 ^ sig_1163;
assign sig_1207 = sig_1159 ^ sig_1158;
assign sig_1224 = A[1] & B[8];
assign sig_1225 = A[1] & B[9];
assign sig_1226 = B[9] & A[0];
assign sig_1227 = A[0] & B[8];
assign sig_1228 = sig_1226 | sig_1224;
assign sig_1229 = A[3] & B[8];
assign sig_1230 = A[3] & B[9];
assign sig_1231 = B[9] & A[2];
assign sig_1232 = A[2] & B[8];
assign sig_1233 = sig_1231 | sig_1229;
assign sig_1234 = A[1] & B[10];
assign sig_1235 = A[1] & B[11];
assign sig_1236 = B[11] & A[0];
assign sig_1237 = A[0] & B[10];
assign sig_1238 = sig_1236 | sig_1234;
assign sig_1239 = A[3] & B[10];
assign sig_1240 = A[3] & B[11];
assign sig_1241 = B[11] & A[2];
assign sig_1242 = A[2] & B[10];
assign sig_1243 = sig_1241 | sig_1239;
assign sig_1248 = sig_1232 ^ sig_1225;
assign sig_1250 = sig_1232 & sig_1225;
assign sig_1255 = sig_1233 & sig_1250;
assign sig_1257 = sig_1230 ^ sig_1242;
assign sig_1258 = sig_1230 & sig_1242;
assign sig_1259 = sig_1257 & sig_1255;
assign sig_1261 = sig_1258 | sig_1259;
assign sig_1263 = sig_1243 & sig_1261;
assign sig_1267 = sig_1240 & sig_1263;
assign sig_1272 = sig_1257 ^ sig_1255;
assign sig_1274 = sig_1240 ^ sig_1263;
assign sig_1275 = sig_1243 ^ sig_1261;
assign sig_1277 = sig_1233 ^ sig_1250;
assign sig_1290 = sig_1237 ^ sig_1248;
assign sig_1292 = sig_1237 & sig_1248;
assign sig_1294 = sig_1238 ^ sig_1277;
assign sig_1296 = sig_1238 & sig_1277;
assign sig_1297 = sig_1294 & sig_1292;
assign sig_1298 = sig_1296 | sig_1297;
assign sig_1299 = sig_1235 ^ sig_1272;
assign sig_1300 = sig_1235 & sig_1272;
assign sig_1301 = sig_1299 & sig_1298;
assign sig_1303 = sig_1300 | sig_1301;
assign sig_1305 = sig_1275 & sig_1303;
assign sig_1309 = sig_1274 & sig_1305;
assign sig_1314 = sig_1299 ^ sig_1298;
assign sig_1315 = sig_1267 ^ sig_1309;
assign sig_1316 = sig_1274 ^ sig_1305;
assign sig_1317 = sig_1275 ^ sig_1303;
assign sig_1319 = sig_1294 ^ sig_1292;
assign sig_1328 = A[5] & B[8];
assign sig_1329 = A[5] & B[9];
assign sig_1330 = B[9] & A[4];
assign sig_1331 = A[4] & B[8];
assign sig_1332 = sig_1330 | sig_1328;
assign sig_1333 = A[7] & B[8];
assign sig_1334 = A[7] & B[9];
assign sig_1335 = B[9] & A[6];
assign sig_1336 = A[6] & B[8];
assign sig_1337 = sig_1335 | sig_1333;
assign sig_1338 = A[5] & B[10];
assign sig_1339 = A[5] & B[11];
assign sig_1340 = B[11] & A[4];
assign sig_1341 = A[4] & B[10];
assign sig_1342 = sig_1340 | sig_1338;
assign sig_1343 = A[7] & B[10];
assign sig_1344 = A[7] & B[11];
assign sig_1345 = B[11] & A[6];
assign sig_1346 = A[6] & B[10];
assign sig_1347 = sig_1345 | sig_1343;
assign sig_1352 = sig_1336 ^ sig_1329;
assign sig_1354 = sig_1336 & sig_1329;
assign sig_1359 = sig_1337 & sig_1354;
assign sig_1361 = sig_1334 ^ sig_1346;
assign sig_1362 = sig_1334 & sig_1346;
assign sig_1363 = sig_1361 & sig_1359;
assign sig_1365 = sig_1362 | sig_1363;
assign sig_1367 = sig_1347 & sig_1365;
assign sig_1371 = sig_1344 & sig_1367;
assign sig_1376 = sig_1361 ^ sig_1359;
assign sig_1378 = sig_1344 ^ sig_1367;
assign sig_1379 = sig_1347 ^ sig_1365;
assign sig_1381 = sig_1337 ^ sig_1354;
assign sig_1394 = sig_1341 ^ sig_1352;
assign sig_1396 = sig_1341 & sig_1352;
assign sig_1398 = sig_1342 ^ sig_1381;
assign sig_1400 = sig_1342 & sig_1381;
assign sig_1401 = sig_1398 & sig_1396;
assign sig_1402 = sig_1400 | sig_1401;
assign sig_1403 = sig_1339 ^ sig_1376;
assign sig_1404 = sig_1339 & sig_1376;
assign sig_1405 = sig_1403 & sig_1402;
assign sig_1407 = sig_1404 | sig_1405;
assign sig_1409 = sig_1379 & sig_1407;
assign sig_1413 = sig_1378 & sig_1409;
assign sig_1418 = sig_1403 ^ sig_1402;
assign sig_1419 = sig_1371 ^ sig_1413;
assign sig_1420 = sig_1378 ^ sig_1409;
assign sig_1421 = sig_1379 ^ sig_1407;
assign sig_1423 = sig_1398 ^ sig_1396;
assign sig_1432 = A[1] & B[12];
assign sig_1433 = A[1] & B[13];
assign sig_1434 = B[13] & A[0];
assign sig_1435 = A[0] & B[12];
assign sig_1436 = sig_1434 | sig_1432;
assign sig_1437 = A[3] & B[12];
assign sig_1438 = A[3] & B[13];
assign sig_1439 = B[13] & A[2];
assign sig_1440 = A[2] & B[12];
assign sig_1441 = sig_1439 | sig_1437;
assign sig_1442 = A[1] & B[14];
assign sig_1443 = A[1] & B[15];
assign sig_1444 = B[15] & A[0];
assign sig_1445 = A[0] & B[14];
assign sig_1446 = sig_1444 | sig_1442;
assign sig_1447 = A[3] & B[14];
assign sig_1448 = A[3] & B[15];
assign sig_1449 = B[15] & A[2];
assign sig_1450 = A[2] & B[14];
assign sig_1451 = sig_1449 | sig_1447;
assign sig_1456 = sig_1440 ^ sig_1433;
assign sig_1458 = sig_1440 & sig_1433;
assign sig_1463 = sig_1441 & sig_1458;
assign sig_1465 = sig_1438 ^ sig_1450;
assign sig_1466 = sig_1438 & sig_1450;
assign sig_1467 = sig_1465 & sig_1463;
assign sig_1469 = sig_1466 | sig_1467;
assign sig_1471 = sig_1451 & sig_1469;
assign sig_1475 = sig_1448 & sig_1471;
assign sig_1480 = sig_1465 ^ sig_1463;
assign sig_1482 = sig_1448 ^ sig_1471;
assign sig_1483 = sig_1451 ^ sig_1469;
assign sig_1485 = sig_1441 ^ sig_1458;
assign sig_1498 = sig_1445 ^ sig_1456;
assign sig_1500 = sig_1445 & sig_1456;
assign sig_1502 = sig_1446 ^ sig_1485;
assign sig_1504 = sig_1446 & sig_1485;
assign sig_1505 = sig_1502 & sig_1500;
assign sig_1506 = sig_1504 | sig_1505;
assign sig_1507 = sig_1443 ^ sig_1480;
assign sig_1508 = sig_1443 & sig_1480;
assign sig_1509 = sig_1507 & sig_1506;
assign sig_1511 = sig_1508 | sig_1509;
assign sig_1513 = sig_1483 & sig_1511;
assign sig_1517 = sig_1482 & sig_1513;
assign sig_1522 = sig_1507 ^ sig_1506;
assign sig_1523 = sig_1475 ^ sig_1517;
assign sig_1524 = sig_1482 ^ sig_1513;
assign sig_1525 = sig_1483 ^ sig_1511;
assign sig_1527 = sig_1502 ^ sig_1500;
assign sig_1536 = A[5] & B[12];
assign sig_1537 = A[5] & B[13];
assign sig_1538 = B[13] & A[4];
assign sig_1539 = A[4] & B[12];
assign sig_1540 = sig_1538 | sig_1536;
assign sig_1541 = A[7] & B[12];
assign sig_1542 = A[7] & B[13];
assign sig_1543 = B[13] & A[6];
assign sig_1544 = A[6] & B[12];
assign sig_1545 = sig_1543 | sig_1541;
assign sig_1546 = A[5] & B[14];
assign sig_1547 = A[5] & B[15];
assign sig_1548 = B[15] & A[4];
assign sig_1549 = A[4] & B[14];
assign sig_1550 = sig_1548 | sig_1546;
assign sig_1551 = A[7] & B[14];
assign sig_1552 = A[7] & B[15];
assign sig_1553 = B[15] & A[6];
assign sig_1554 = A[6] & B[14];
assign sig_1555 = sig_1553 | sig_1551;
assign sig_1560 = sig_1544 ^ sig_1537;
assign sig_1562 = sig_1544 & sig_1537;
assign sig_1567 = sig_1545 & sig_1562;
assign sig_1569 = sig_1542 ^ sig_1554;
assign sig_1570 = sig_1542 & sig_1554;
assign sig_1571 = sig_1569 & sig_1567;
assign sig_1573 = sig_1570 | sig_1571;
assign sig_1575 = sig_1555 & sig_1573;
assign sig_1579 = sig_1552 & sig_1575;
assign sig_1584 = sig_1569 ^ sig_1567;
assign sig_1586 = sig_1552 ^ sig_1575;
assign sig_1587 = sig_1555 ^ sig_1573;
assign sig_1589 = sig_1545 ^ sig_1562;
assign sig_1602 = sig_1549 ^ sig_1560;
assign sig_1604 = sig_1549 & sig_1560;
assign sig_1606 = sig_1550 ^ sig_1589;
assign sig_1608 = sig_1550 & sig_1589;
assign sig_1609 = sig_1606 & sig_1604;
assign sig_1610 = sig_1608 | sig_1609;
assign sig_1611 = sig_1547 ^ sig_1584;
assign sig_1612 = sig_1547 & sig_1584;
assign sig_1613 = sig_1611 & sig_1610;
assign sig_1615 = sig_1612 | sig_1613;
assign sig_1617 = sig_1587 & sig_1615;
assign sig_1621 = sig_1586 & sig_1617;
assign sig_1626 = sig_1611 ^ sig_1610;
assign sig_1627 = sig_1579 ^ sig_1621;
assign sig_1628 = sig_1586 ^ sig_1617;
assign sig_1629 = sig_1587 ^ sig_1615;
assign sig_1631 = sig_1606 ^ sig_1604;
assign sig_1652 = sig_1331 ^ sig_1314;
assign sig_1654 = sig_1331 & sig_1314;
assign sig_1656 = sig_1332 ^ sig_1317;
assign sig_1658 = sig_1656 & sig_1654;
assign sig_1659 = sig_1332 & sig_1317;
assign sig_1660 = sig_1659 | sig_1658;
assign sig_1661 = sig_1394 ^ sig_1316;
assign sig_1662 = sig_1661 & sig_1660;
assign sig_1663 = sig_1394 & sig_1316;
assign sig_1664 = sig_1663 | sig_1662;
assign sig_1665 = sig_1423 ^ sig_1315;
assign sig_1666 = sig_1665 & sig_1664;
assign sig_1667 = sig_1423 & sig_1315;
assign sig_1668 = sig_1418 ^ sig_1539;
assign sig_1669 = sig_1667 | sig_1666;
assign sig_1670 = sig_1418 & sig_1539;
assign sig_1671 = sig_1668 & sig_1669;
assign sig_1672 = sig_1421 ^ sig_1540;
assign sig_1673 = sig_1670 | sig_1671;
assign sig_1674 = sig_1421 & sig_1540;
assign sig_1675 = sig_1672 & sig_1673;
assign sig_1676 = sig_1420 ^ sig_1602;
assign sig_1677 = sig_1674 | sig_1675;
assign sig_1678 = sig_1676 & sig_1677;
assign sig_1679 = sig_1420 & sig_1602;
assign sig_1680 = sig_1679 | sig_1678;
assign sig_1681 = sig_1419 ^ sig_1631;
assign sig_1682 = sig_1681 & sig_1680;
assign sig_1683 = sig_1419 & sig_1631;
assign sig_1684 = sig_1683 | sig_1682;
assign sig_1686 = sig_1626 & sig_1684;
assign sig_1691 = sig_1629 & sig_1686;
assign sig_1694 = sig_1628 & sig_1691;
assign sig_1698 = sig_1656 ^ sig_1654;
assign sig_1701 = sig_1676 ^ sig_1677;
assign sig_1702 = sig_1661 ^ sig_1660;
assign sig_1703 = sig_1681 ^ sig_1680;
assign sig_1704 = sig_1626 ^ sig_1684;
assign sig_1707 = sig_1629 ^ sig_1686;
assign sig_1708 = sig_1628 ^ sig_1691;
assign sig_1709 = sig_1672 ^ sig_1673;
assign sig_1711 = sig_1627 ^ sig_1694;
assign sig_1712 = sig_1668 ^ sig_1669;
assign sig_1713 = sig_1665 ^ sig_1664;
assign sig_1742 = sig_1435 ^ sig_1652;
assign sig_1744 = sig_1435 & sig_1652;
assign sig_1746 = sig_1436 ^ sig_1698;
assign sig_1748 = sig_1746 & sig_1744;
assign sig_1749 = sig_1436 & sig_1698;
assign sig_1750 = sig_1749 | sig_1748;
assign sig_1751 = sig_1498 ^ sig_1702;
assign sig_1752 = sig_1751 & sig_1750;
assign sig_1753 = sig_1498 & sig_1702;
assign sig_1754 = sig_1753 | sig_1752;
assign sig_1755 = sig_1527 ^ sig_1713;
assign sig_1756 = sig_1755 & sig_1754;
assign sig_1757 = sig_1527 & sig_1713;
assign sig_1758 = sig_1522 ^ sig_1712;
assign sig_1759 = sig_1757 | sig_1756;
assign sig_1760 = sig_1522 & sig_1712;
assign sig_1761 = sig_1758 & sig_1759;
assign sig_1762 = sig_1525 ^ sig_1709;
assign sig_1763 = sig_1760 | sig_1761;
assign sig_1764 = sig_1525 & sig_1709;
assign sig_1765 = sig_1762 & sig_1763;
assign sig_1766 = sig_1524 ^ sig_1701;
assign sig_1767 = sig_1764 | sig_1765;
assign sig_1768 = sig_1766 & sig_1767;
assign sig_1769 = sig_1524 & sig_1701;
assign sig_1770 = sig_1769 | sig_1768;
assign sig_1771 = sig_1523 ^ sig_1703;
assign sig_1772 = sig_1771 & sig_1770;
assign sig_1773 = sig_1523 & sig_1703;
assign sig_1774 = sig_1773 | sig_1772;
assign sig_1776 = sig_1704 & sig_1774;
assign sig_1781 = sig_1707 & sig_1776;
assign sig_1784 = sig_1708 & sig_1781;
assign sig_1788 = sig_1746 ^ sig_1744;
assign sig_1791 = sig_1766 ^ sig_1767;
assign sig_1792 = sig_1751 ^ sig_1750;
assign sig_1793 = sig_1771 ^ sig_1770;
assign sig_1794 = sig_1704 ^ sig_1774;
assign sig_1797 = sig_1707 ^ sig_1776;
assign sig_1798 = sig_1708 ^ sig_1781;
assign sig_1799 = sig_1762 ^ sig_1763;
assign sig_1801 = sig_1711 ^ sig_1784;
assign sig_1802 = sig_1758 ^ sig_1759;
assign sig_1803 = sig_1755 ^ sig_1754;
assign sig_1820 = A[9] & B[8];
assign sig_1821 = A[9] & B[9];
assign sig_1822 = B[9] & A[8];
assign sig_1823 = A[8] & B[8];
assign sig_1824 = sig_1822 | sig_1820;
assign sig_1825 = A[11] & B[8];
assign sig_1826 = A[11] & B[9];
assign sig_1827 = B[9] & A[10];
assign sig_1828 = A[10] & B[8];
assign sig_1829 = sig_1827 | sig_1825;
assign sig_1830 = A[9] & B[10];
assign sig_1831 = A[9] & B[11];
assign sig_1832 = B[11] & A[8];
assign sig_1833 = A[8] & B[10];
assign sig_1834 = sig_1832 | sig_1830;
assign sig_1835 = A[11] & B[10];
assign sig_1836 = A[11] & B[11];
assign sig_1837 = B[11] & A[10];
assign sig_1838 = A[10] & B[10];
assign sig_1839 = sig_1837 | sig_1835;
assign sig_1844 = sig_1828 ^ sig_1821;
assign sig_1846 = sig_1828 & sig_1821;
assign sig_1851 = sig_1829 & sig_1846;
assign sig_1853 = sig_1826 ^ sig_1838;
assign sig_1854 = sig_1826 & sig_1838;
assign sig_1855 = sig_1853 & sig_1851;
assign sig_1857 = sig_1854 | sig_1855;
assign sig_1859 = sig_1839 & sig_1857;
assign sig_1863 = sig_1836 & sig_1859;
assign sig_1868 = sig_1853 ^ sig_1851;
assign sig_1870 = sig_1836 ^ sig_1859;
assign sig_1871 = sig_1839 ^ sig_1857;
assign sig_1873 = sig_1829 ^ sig_1846;
assign sig_1886 = sig_1833 ^ sig_1844;
assign sig_1888 = sig_1833 & sig_1844;
assign sig_1890 = sig_1834 ^ sig_1873;
assign sig_1892 = sig_1834 & sig_1873;
assign sig_1893 = sig_1890 & sig_1888;
assign sig_1894 = sig_1892 | sig_1893;
assign sig_1895 = sig_1831 ^ sig_1868;
assign sig_1896 = sig_1831 & sig_1868;
assign sig_1897 = sig_1895 & sig_1894;
assign sig_1899 = sig_1896 | sig_1897;
assign sig_1901 = sig_1871 & sig_1899;
assign sig_1905 = sig_1870 & sig_1901;
assign sig_1910 = sig_1895 ^ sig_1894;
assign sig_1911 = sig_1863 ^ sig_1905;
assign sig_1912 = sig_1870 ^ sig_1901;
assign sig_1913 = sig_1871 ^ sig_1899;
assign sig_1915 = sig_1890 ^ sig_1888;
assign sig_1924 = A[13] & B[8];
assign sig_1925 = A[13] & B[9];
assign sig_1926 = B[9] & A[12];
assign sig_1927 = A[12] & B[8];
assign sig_1928 = sig_1926 | sig_1924;
assign sig_1929 = A[15] & B[8];
assign sig_1930 = A[15] & B[9];
assign sig_1931 = B[9] & A[14];
assign sig_1932 = A[14] & B[8];
assign sig_1933 = sig_1931 | sig_1929;
assign sig_1934 = A[13] & B[10];
assign sig_1935 = A[13] & B[11];
assign sig_1936 = B[11] & A[12];
assign sig_1937 = A[12] & B[10];
assign sig_1938 = sig_1936 | sig_1934;
assign sig_1939 = A[15] & B[10];
assign sig_1940 = A[15] & B[11];
assign sig_1941 = B[11] & A[14];
assign sig_1942 = A[14] & B[10];
assign sig_1943 = sig_1941 | sig_1939;
assign sig_1948 = sig_1932 ^ sig_1925;
assign sig_1950 = sig_1932 & sig_1925;
assign sig_1955 = sig_1933 & sig_1950;
assign sig_1957 = sig_1930 ^ sig_1942;
assign sig_1958 = sig_1930 & sig_1942;
assign sig_1959 = sig_1957 & sig_1955;
assign sig_1961 = sig_1958 | sig_1959;
assign sig_1963 = sig_1943 & sig_1961;
assign sig_1967 = sig_1940 & sig_1963;
assign sig_1972 = sig_1957 ^ sig_1955;
assign sig_1974 = sig_1940 ^ sig_1963;
assign sig_1975 = sig_1943 ^ sig_1961;
assign sig_1977 = sig_1933 ^ sig_1950;
assign sig_1990 = sig_1937 ^ sig_1948;
assign sig_1992 = sig_1937 & sig_1948;
assign sig_1994 = sig_1938 ^ sig_1977;
assign sig_1996 = sig_1938 & sig_1977;
assign sig_1997 = sig_1994 & sig_1992;
assign sig_1998 = sig_1996 | sig_1997;
assign sig_1999 = sig_1935 ^ sig_1972;
assign sig_2000 = sig_1935 & sig_1972;
assign sig_2001 = sig_1999 & sig_1998;
assign sig_2003 = sig_2000 | sig_2001;
assign sig_2005 = sig_1975 & sig_2003;
assign sig_2009 = sig_1974 & sig_2005;
assign sig_2014 = sig_1999 ^ sig_1998;
assign sig_2015 = sig_1967 ^ sig_2009;
assign sig_2016 = sig_1974 ^ sig_2005;
assign sig_2017 = sig_1975 ^ sig_2003;
assign sig_2019 = sig_1994 ^ sig_1992;
assign sig_2028 = A[9] & B[12];
assign sig_2029 = A[9] & B[13];
assign sig_2030 = B[13] & A[8];
assign sig_2031 = A[8] & B[12];
assign sig_2032 = sig_2030 | sig_2028;
assign sig_2033 = A[11] & B[12];
assign sig_2034 = A[11] & B[13];
assign sig_2035 = B[13] & A[10];
assign sig_2036 = A[10] & B[12];
assign sig_2037 = sig_2035 | sig_2033;
assign sig_2038 = A[9] & B[14];
assign sig_2039 = A[9] & B[15];
assign sig_2040 = B[15] & A[8];
assign sig_2041 = A[8] & B[14];
assign sig_2042 = sig_2040 | sig_2038;
assign sig_2043 = A[11] & B[14];
assign sig_2044 = A[11] & B[15];
assign sig_2045 = B[15] & A[10];
assign sig_2046 = A[10] & B[14];
assign sig_2047 = sig_2045 | sig_2043;
assign sig_2052 = sig_2036 ^ sig_2029;
assign sig_2054 = sig_2036 & sig_2029;
assign sig_2059 = sig_2037 & sig_2054;
assign sig_2061 = sig_2034 ^ sig_2046;
assign sig_2062 = sig_2034 & sig_2046;
assign sig_2063 = sig_2061 & sig_2059;
assign sig_2065 = sig_2062 | sig_2063;
assign sig_2067 = sig_2047 & sig_2065;
assign sig_2071 = sig_2044 & sig_2067;
assign sig_2076 = sig_2061 ^ sig_2059;
assign sig_2078 = sig_2044 ^ sig_2067;
assign sig_2079 = sig_2047 ^ sig_2065;
assign sig_2081 = sig_2037 ^ sig_2054;
assign sig_2094 = sig_2041 ^ sig_2052;
assign sig_2096 = sig_2041 & sig_2052;
assign sig_2098 = sig_2042 ^ sig_2081;
assign sig_2100 = sig_2042 & sig_2081;
assign sig_2101 = sig_2098 & sig_2096;
assign sig_2102 = sig_2100 | sig_2101;
assign sig_2103 = sig_2039 ^ sig_2076;
assign sig_2104 = sig_2039 & sig_2076;
assign sig_2105 = sig_2103 & sig_2102;
assign sig_2107 = sig_2104 | sig_2105;
assign sig_2109 = sig_2079 & sig_2107;
assign sig_2113 = sig_2078 & sig_2109;
assign sig_2118 = sig_2103 ^ sig_2102;
assign sig_2119 = sig_2071 ^ sig_2113;
assign sig_2120 = sig_2078 ^ sig_2109;
assign sig_2121 = sig_2079 ^ sig_2107;
assign sig_2123 = sig_2098 ^ sig_2096;
assign sig_2132 = A[13] & B[12];
assign sig_2133 = A[13] & B[13];
assign sig_2134 = B[13] & A[12];
assign sig_2135 = A[12] & B[12];
assign sig_2136 = sig_2134 | sig_2132;
assign sig_2137 = A[15] & B[12];
assign sig_2138 = A[15] & B[13];
assign sig_2139 = B[13] & A[14];
assign sig_2140 = A[14] & B[12];
assign sig_2141 = sig_2139 | sig_2137;
assign sig_2142 = A[13] & B[14];
assign sig_2143 = A[13] & B[15];
assign sig_2144 = B[15] & A[12];
assign sig_2145 = A[12] & B[14];
assign sig_2146 = sig_2144 | sig_2142;
assign sig_2147 = A[15] & B[14];
assign sig_2148 = A[15] & B[15];
assign sig_2149 = B[15] & A[14];
assign sig_2150 = A[14] & B[14];
assign sig_2151 = sig_2149 | sig_2147;
assign sig_2156 = sig_2140 ^ sig_2133;
assign sig_2158 = sig_2140 & sig_2133;
assign sig_2163 = sig_2141 & sig_2158;
assign sig_2165 = sig_2138 ^ sig_2150;
assign sig_2166 = sig_2138 & sig_2150;
assign sig_2167 = sig_2165 & sig_2163;
assign sig_2169 = sig_2166 | sig_2167;
assign sig_2171 = sig_2151 & sig_2169;
assign sig_2175 = sig_2148 & sig_2171;
assign sig_2180 = sig_2165 ^ sig_2163;
assign sig_2182 = sig_2148 ^ sig_2171;
assign sig_2183 = sig_2151 ^ sig_2169;
assign sig_2185 = sig_2141 ^ sig_2158;
assign sig_2198 = sig_2145 ^ sig_2156;
assign sig_2200 = sig_2145 & sig_2156;
assign sig_2202 = sig_2146 ^ sig_2185;
assign sig_2204 = sig_2146 & sig_2185;
assign sig_2205 = sig_2202 & sig_2200;
assign sig_2206 = sig_2204 | sig_2205;
assign sig_2207 = sig_2143 ^ sig_2180;
assign sig_2208 = sig_2143 & sig_2180;
assign sig_2209 = sig_2207 & sig_2206;
assign sig_2211 = sig_2208 | sig_2209;
assign sig_2213 = sig_2183 & sig_2211;
assign sig_2217 = sig_2182 & sig_2213;
assign sig_2222 = sig_2207 ^ sig_2206;
assign sig_2223 = sig_2175 ^ sig_2217;
assign sig_2224 = sig_2182 ^ sig_2213;
assign sig_2225 = sig_2183 ^ sig_2211;
assign sig_2227 = sig_2202 ^ sig_2200;
assign sig_2248 = sig_1927 ^ sig_1910;
assign sig_2250 = sig_1927 & sig_1910;
assign sig_2252 = sig_1928 ^ sig_1913;
assign sig_2254 = sig_2252 & sig_2250;
assign sig_2255 = sig_1928 & sig_1913;
assign sig_2256 = sig_2255 | sig_2254;
assign sig_2257 = sig_1990 ^ sig_1912;
assign sig_2258 = sig_2257 & sig_2256;
assign sig_2259 = sig_1990 & sig_1912;
assign sig_2260 = sig_2259 | sig_2258;
assign sig_2261 = sig_2019 ^ sig_1911;
assign sig_2262 = sig_2261 & sig_2260;
assign sig_2263 = sig_2019 & sig_1911;
assign sig_2264 = sig_2014 ^ sig_2135;
assign sig_2265 = sig_2263 | sig_2262;
assign sig_2266 = sig_2014 & sig_2135;
assign sig_2267 = sig_2264 & sig_2265;
assign sig_2268 = sig_2017 ^ sig_2136;
assign sig_2269 = sig_2266 | sig_2267;
assign sig_2270 = sig_2017 & sig_2136;
assign sig_2271 = sig_2268 & sig_2269;
assign sig_2272 = sig_2016 ^ sig_2198;
assign sig_2273 = sig_2270 | sig_2271;
assign sig_2274 = sig_2272 & sig_2273;
assign sig_2275 = sig_2016 & sig_2198;
assign sig_2276 = sig_2275 | sig_2274;
assign sig_2277 = sig_2015 ^ sig_2227;
assign sig_2278 = sig_2277 & sig_2276;
assign sig_2279 = sig_2015 & sig_2227;
assign sig_2280 = sig_2279 | sig_2278;
assign sig_2282 = sig_2222 & sig_2280;
assign sig_2287 = sig_2225 & sig_2282;
assign sig_2290 = sig_2224 & sig_2287;
assign sig_2294 = sig_2252 ^ sig_2250;
assign sig_2297 = sig_2272 ^ sig_2273;
assign sig_2298 = sig_2257 ^ sig_2256;
assign sig_2299 = sig_2277 ^ sig_2276;
assign sig_2300 = sig_2222 ^ sig_2280;
assign sig_2303 = sig_2225 ^ sig_2282;
assign sig_2304 = sig_2224 ^ sig_2287;
assign sig_2305 = sig_2268 ^ sig_2269;
assign sig_2307 = sig_2223 ^ sig_2290;
assign sig_2308 = sig_2264 ^ sig_2265;
assign sig_2309 = sig_2261 ^ sig_2260;
assign sig_2338 = sig_2031 ^ sig_2248;
assign sig_2340 = sig_2031 & sig_2248;
assign sig_2342 = sig_2032 ^ sig_2294;
assign sig_2344 = sig_2342 & sig_2340;
assign sig_2345 = sig_2032 & sig_2294;
assign sig_2346 = sig_2345 | sig_2344;
assign sig_2347 = sig_2094 ^ sig_2298;
assign sig_2348 = sig_2347 & sig_2346;
assign sig_2349 = sig_2094 & sig_2298;
assign sig_2350 = sig_2349 | sig_2348;
assign sig_2351 = sig_2123 ^ sig_2309;
assign sig_2352 = sig_2351 & sig_2350;
assign sig_2353 = sig_2123 & sig_2309;
assign sig_2354 = sig_2118 ^ sig_2308;
assign sig_2355 = sig_2353 | sig_2352;
assign sig_2356 = sig_2118 & sig_2308;
assign sig_2357 = sig_2354 & sig_2355;
assign sig_2358 = sig_2121 ^ sig_2305;
assign sig_2359 = sig_2356 | sig_2357;
assign sig_2360 = sig_2121 & sig_2305;
assign sig_2361 = sig_2358 & sig_2359;
assign sig_2362 = sig_2120 ^ sig_2297;
assign sig_2363 = sig_2360 | sig_2361;
assign sig_2364 = sig_2362 & sig_2363;
assign sig_2365 = sig_2120 & sig_2297;
assign sig_2366 = sig_2365 | sig_2364;
assign sig_2367 = sig_2119 ^ sig_2299;
assign sig_2368 = sig_2367 & sig_2366;
assign sig_2369 = sig_2119 & sig_2299;
assign sig_2370 = sig_2369 | sig_2368;
assign sig_2372 = sig_2300 & sig_2370;
assign sig_2377 = sig_2303 & sig_2372;
assign sig_2380 = sig_2304 & sig_2377;
assign sig_2384 = sig_2342 ^ sig_2340;
assign sig_2387 = sig_2362 ^ sig_2363;
assign sig_2388 = sig_2347 ^ sig_2346;
assign sig_2389 = sig_2367 ^ sig_2366;
assign sig_2390 = sig_2300 ^ sig_2370;
assign sig_2393 = sig_2303 ^ sig_2372;
assign sig_2394 = sig_2304 ^ sig_2377;
assign sig_2395 = sig_2358 ^ sig_2359;
assign sig_2397 = sig_2307 ^ sig_2380;
assign sig_2398 = sig_2354 ^ sig_2355;
assign sig_2399 = sig_2351 ^ sig_2350;
assign sig_2432 = sig_631 ^ sig_610;
assign sig_2433 = sig_631 & sig_610;
assign sig_2434 = sig_632 ^ sig_607;
assign sig_2435 = sig_632 & sig_607;
assign sig_2436 = sig_694 ^ sig_599;
assign sig_2437 = sig_694 & sig_599;
assign sig_2438 = sig_723 ^ sig_601;
assign sig_2439 = sig_723 & sig_601;
assign sig_2440 = sig_1146 ^ sig_602;
assign sig_2441 = sig_1146 & sig_602;
assign sig_2442 = sig_1192 ^ sig_605;
assign sig_2443 = sig_1192 & sig_605;
assign sig_2444 = sig_1196 ^ sig_606;
assign sig_2445 = sig_1196 & sig_606;
assign sig_2446 = sig_1207 ^ sig_609;
assign sig_2447 = sig_1207 & sig_609;
assign sig_2448 = sig_1206 ^ sig_1823;
assign sig_2449 = sig_1206 & sig_1823;
assign sig_2450 = sig_1203 ^ sig_1824;
assign sig_2451 = sig_1203 & sig_1824;
assign sig_2452 = sig_1195 ^ sig_1886;
assign sig_2453 = sig_1195 & sig_1886;
assign sig_2454 = sig_1197 ^ sig_1915;
assign sig_2455 = sig_1197 & sig_1915;
assign sig_2456 = sig_1198 ^ sig_2338;
assign sig_2457 = sig_1198 & sig_2338;
assign sig_2458 = sig_1201 ^ sig_2384;
assign sig_2459 = sig_1201 & sig_2384;
assign sig_2460 = sig_1202 ^ sig_2388;
assign sig_2461 = sig_1202 & sig_2388;
assign sig_2462 = sig_1205 ^ sig_2399;
assign sig_2463 = sig_1205 & sig_2399;
assign sig_2503 = sig_2434 ^ sig_2433;
assign sig_2504 = sig_2434 & sig_2433;
assign sig_2505 = sig_2435 | sig_2504;
assign sig_2506 = sig_2436 ^ sig_2505;
assign sig_2507 = sig_2436 & sig_2505;
assign sig_2508 = sig_2437 | sig_2507;
assign sig_2509 = sig_2438 ^ sig_2508;
assign sig_2510 = sig_2438 & sig_2508;
assign sig_2511 = sig_2439 | sig_2510;
assign sig_2512 = sig_2440 ^ sig_2511;
assign sig_2513 = sig_2440 & sig_2511;
assign sig_2514 = sig_2441 | sig_2513;
assign sig_2515 = sig_2442 ^ sig_2514;
assign sig_2516 = sig_2442 & sig_2514;
assign sig_2517 = sig_2443 | sig_2516;
assign sig_2518 = sig_2444 ^ sig_2517;
assign sig_2519 = sig_2444 & sig_2517;
assign sig_2520 = sig_2445 | sig_2519;
assign sig_2521 = sig_2446 ^ sig_2520;
assign sig_2522 = sig_2446 & sig_2520;
assign sig_2523 = sig_2447 | sig_2522;
assign sig_2524 = sig_2448 ^ sig_2523;
assign sig_2525 = sig_2448 & sig_2523;
assign sig_2526 = sig_2449 | sig_2525;
assign sig_2527 = sig_2450 ^ sig_2526;
assign sig_2528 = sig_2450 & sig_2526;
assign sig_2529 = sig_2451 | sig_2528;
assign sig_2530 = sig_2452 ^ sig_2529;
assign sig_2531 = sig_2452 & sig_2529;
assign sig_2532 = sig_2453 | sig_2531;
assign sig_2533 = sig_2454 ^ sig_2532;
assign sig_2534 = sig_2454 & sig_2532;
assign sig_2535 = sig_2455 | sig_2534;
assign sig_2536 = sig_2456 ^ sig_2535;
assign sig_2537 = sig_2456 & sig_2535;
assign sig_2538 = sig_2457 | sig_2537;
assign sig_2539 = sig_2458 ^ sig_2538;
assign sig_2540 = sig_2458 & sig_2538;
assign sig_2541 = sig_2459 | sig_2540;
assign sig_2542 = sig_2460 ^ sig_2541;
assign sig_2543 = sig_2460 & sig_2541;
assign sig_2544 = sig_2461 | sig_2543;
assign sig_2545 = sig_2462 ^ sig_2544;
assign sig_2546 = sig_2462 & sig_2544;
assign sig_2547 = sig_2463 | sig_2546;
assign sig_2548 = sig_2398 ^ sig_2547;
assign sig_2549 = sig_2398 & sig_2547;
assign sig_2551 = sig_2395 ^ sig_2549;
assign sig_2552 = sig_2395 & sig_2549;
assign sig_2554 = sig_2387 ^ sig_2552;
assign sig_2555 = sig_2387 & sig_2552;
assign sig_2557 = sig_2389 ^ sig_2555;
assign sig_2558 = sig_2389 & sig_2555;
assign sig_2560 = sig_2390 ^ sig_2558;
assign sig_2561 = sig_2390 & sig_2558;
assign sig_2563 = sig_2393 ^ sig_2561;
assign sig_2564 = sig_2393 & sig_2561;
assign sig_2566 = sig_2394 ^ sig_2564;
assign sig_2567 = sig_2394 & sig_2564;
assign sig_2569 = sig_2397 ^ sig_2567;
assign sig_2586 = sig_1227 ^ sig_2432;
assign sig_2587 = sig_1227 & sig_2432;
assign sig_2588 = sig_1228 ^ sig_2503;
assign sig_2589 = sig_1228 & sig_2503;
assign sig_2590 = sig_1290 ^ sig_2506;
assign sig_2591 = sig_1290 & sig_2506;
assign sig_2592 = sig_1319 ^ sig_2509;
assign sig_2593 = sig_1319 & sig_2509;
assign sig_2594 = sig_1742 ^ sig_2512;
assign sig_2595 = sig_1742 & sig_2512;
assign sig_2596 = sig_1788 ^ sig_2515;
assign sig_2597 = sig_1788 & sig_2515;
assign sig_2598 = sig_1792 ^ sig_2518;
assign sig_2599 = sig_1792 & sig_2518;
assign sig_2600 = sig_1803 ^ sig_2521;
assign sig_2601 = sig_1803 & sig_2521;
assign sig_2602 = sig_1802 ^ sig_2524;
assign sig_2603 = sig_1802 & sig_2524;
assign sig_2604 = sig_1799 ^ sig_2527;
assign sig_2605 = sig_1799 & sig_2527;
assign sig_2606 = sig_1791 ^ sig_2530;
assign sig_2607 = sig_1791 & sig_2530;
assign sig_2608 = sig_1793 ^ sig_2533;
assign sig_2609 = sig_1793 & sig_2533;
assign sig_2610 = sig_1794 ^ sig_2536;
assign sig_2611 = sig_1794 & sig_2536;
assign sig_2612 = sig_1797 ^ sig_2539;
assign sig_2613 = sig_1797 & sig_2539;
assign sig_2614 = sig_1798 ^ sig_2542;
assign sig_2615 = sig_1798 & sig_2542;
assign sig_2616 = sig_1801 ^ sig_2545;
assign sig_2617 = sig_1801 & sig_2545;
assign sig_2657 = sig_2588 ^ sig_2587;
assign sig_2658 = sig_2588 & sig_2587;
assign sig_2659 = sig_2589 | sig_2658;
assign sig_2660 = sig_2590 ^ sig_2659;
assign sig_2661 = sig_2590 & sig_2659;
assign sig_2662 = sig_2591 | sig_2661;
assign sig_2663 = sig_2592 ^ sig_2662;
assign sig_2664 = sig_2592 & sig_2662;
assign sig_2665 = sig_2593 | sig_2664;
assign sig_2666 = sig_2594 ^ sig_2665;
assign sig_2667 = sig_2594 & sig_2665;
assign sig_2668 = sig_2595 | sig_2667;
assign sig_2669 = sig_2596 ^ sig_2668;
assign sig_2670 = sig_2596 & sig_2668;
assign sig_2671 = sig_2597 | sig_2670;
assign sig_2672 = sig_2598 ^ sig_2671;
assign sig_2673 = sig_2598 & sig_2671;
assign sig_2674 = sig_2599 | sig_2673;
assign sig_2675 = sig_2600 ^ sig_2674;
assign sig_2676 = sig_2600 & sig_2674;
assign sig_2677 = sig_2601 | sig_2676;
assign sig_2678 = sig_2602 ^ sig_2677;
assign sig_2679 = sig_2602 & sig_2677;
assign sig_2680 = sig_2603 | sig_2679;
assign sig_2681 = sig_2604 ^ sig_2680;
assign sig_2682 = sig_2604 & sig_2680;
assign sig_2683 = sig_2605 | sig_2682;
assign sig_2684 = sig_2606 ^ sig_2683;
assign sig_2685 = sig_2606 & sig_2683;
assign sig_2686 = sig_2607 | sig_2685;
assign sig_2687 = sig_2608 ^ sig_2686;
assign sig_2688 = sig_2608 & sig_2686;
assign sig_2689 = sig_2609 | sig_2688;
assign sig_2690 = sig_2610 ^ sig_2689;
assign sig_2691 = sig_2610 & sig_2689;
assign sig_2692 = sig_2611 | sig_2691;
assign sig_2693 = sig_2612 ^ sig_2692;
assign sig_2694 = sig_2612 & sig_2692;
assign sig_2695 = sig_2613 | sig_2694;
assign sig_2696 = sig_2614 ^ sig_2695;
assign sig_2697 = sig_2614 & sig_2695;
assign sig_2698 = sig_2615 | sig_2697;
assign sig_2699 = sig_2616 ^ sig_2698;
assign sig_2700 = sig_2616 & sig_2698;
assign sig_2701 = sig_2617 | sig_2700;
assign sig_2702 = sig_2548 ^ sig_2701;
assign sig_2703 = sig_2548 & sig_2701;
assign sig_2705 = sig_2551 ^ sig_2703;
assign sig_2706 = sig_2551 & sig_2703;
assign sig_2708 = sig_2554 ^ sig_2706;
assign sig_2709 = sig_2554 & sig_2706;
assign sig_2711 = sig_2557 ^ sig_2709;
assign sig_2712 = sig_2557 & sig_2709;
assign sig_2714 = sig_2560 ^ sig_2712;
assign sig_2715 = sig_2560 & sig_2712;
assign sig_2717 = sig_2563 ^ sig_2715;
assign sig_2718 = sig_2563 & sig_2715;
assign sig_2720 = sig_2566 ^ sig_2718;
assign sig_2721 = sig_2566 & sig_2718;
assign sig_2723 = sig_2569 ^ sig_2721;

assign O[31] = sig_2723;
assign O[30] = sig_2720;
assign O[29] = sig_2717;
assign O[28] = sig_2714;
assign O[27] = sig_2711;
assign O[26] = sig_2708;
assign O[25] = sig_2705;
assign O[24] = sig_2702;
assign O[23] = sig_2699;
assign O[22] = sig_2696;
assign O[21] = sig_2693;
assign O[20] = sig_2690;
assign O[19] = sig_2687;
assign O[18] = sig_2684;
assign O[17] = sig_2681;
assign O[16] = sig_2678;
assign O[15] = sig_2675;
assign O[14] = sig_2672;
assign O[13] = sig_2669;
assign O[12] = sig_2666;
assign O[11] = sig_2663;
assign O[10] = sig_2660;
assign O[9] = sig_2657;
assign O[8] = sig_2586;
assign O[7] = sig_611;
assign O[6] = sig_600;
assign O[5] = sig_596;
assign O[4] = sig_550;
assign O[3] = sig_127;
assign O[2] = sig_98;
assign O[1] = sig_36;
assign O[0] = sig_35;

endmodule


