/***
    * This code is a part of ApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under a XXXX public license.
    * When used, please cite the following article: tbd 
    * This file is pareto optimal sub-set in the pwr and wce parameters
    ***/
    
module mul12u_pwr_0_680_wce_00_0493(A, B, O);
  input [11:0] A, B;
  output [23:0] O;
  wire n_1192, n_1750, n_1751, n_1206, n_1759, n_1613, n_1612, n_1200, n_1816, n_1684;
  wire n_322, n_1105, n_1104, n_1295, n_1294, n_150, n_1866, n_230, n_1758, n_2032;
  wire n_2033, n_126, n_1032, n_428, n_429, n_1402, n_1403, n_1969, n_1968, n_18;
  wire n_19, n_16, n_17, n_1961, n_15, n_12, n_13, n_10, n_11, n_880;
  wire n_1532, n_1714, n_1243, n_1084, n_1085, n_1496, n_1322, n_1916, n_1917, n_1910;
  wire n_1911, n_938, n_1148, n_1662, n_1394, n_1395, n_1983, n_1982, n_1822, n_286;
  wire n_287, n_518, n_794, n_604, n_605, n_795, n_764, n_1932, n_947, n_946;
  wire n_417, n_416, n_1947, n_1366, n_1946, n_45, n_44, n_47, n_46, n_41;
  wire n_40, n_43, n_42, n_1040, n_866, n_1591, n_1895, n_1894, n_460, n_461;
  wire n_1563, n_1562, n_1446, n_1447, n_453, n_1569, n_1568, n_1626, n_1627, n_1620;
  wire n_1621, n_1184, n_1214, n_1743, n_1742, n_1692, n_1874, n_228, n_229, n_185;
  wire n_184, n_2027, n_2026, n_526, n_136, n_137, n_1004, n_1554, n_1555, n_1526;
  wire n_1251, n_1250, n_1700, n_1706, n_1259, n_1258, n_1858, n_1091, n_1090, n_852;
  wire n_1099, n_1098, n_858, n_1316, n_78, n_76, n_77, n_70, n_71, n_1903;
  wire n_1902, n_1417, n_1416, n_1598, n_1411, n_1410, n_1794, n_1795, n_1170, n_1178;
  wire n_1599, n_1772, n_1773, n_1678, n_1778, n_1779, n_1380, n_1830, n_1836, n_917;
  wire n_706, n_700, n_916, n_380, n_2018, n_2019, n_388, n_2010, n_2011, n_778;
  wire n_779, n_772, n_773, n_952, n_953, n_1358, n_1424, n_1425, n_1352, n_30;
  wire n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_1585;
  wire n_1584, n_1048, n_1590, n_1953, n_787, n_1510, n_786, n_1952, n_1453, n_1452;
  wire n_1518, n_1634, n_925, n_924, n_1736, n_1737, n_64, n_1642, n_1127, n_1126;
  wire n_1121, n_1120, n_1844, n_626, n_627, n_620, n_621, n_14, n_1960, n_452;
  wire n_532, n_1648, n_105, n_104, n_1018, n_366, n_1010, n_1540, n_692, n_2041;
  wire n_2040, n_214, n_1264, n_1265, n_1308, n_961, n_960, n_1938, n_1939, n_66;
  wire n_65, n_1933, n_63, n_62, n_1460, n_1461, n_1468, n_1670, n_1787, n_1786;
  wire n_1162, n_8, n_9, n_4, n_5, n_6, n_7, n_0, n_1, n_2;
  wire n_3, n_1765, n_1764, n_1604, n_1605, n_1800, n_1808, n_1242, n_548, n_540;
  wire n_1112, n_1113, n_1286, n_1287, n_714, n_2005, n_2004, n_1026, n_1438, n_1433;
  wire n_1432, n_23, n_22, n_21, n_20, n_27, n_26, n_25, n_24, n_1974;
  wire n_1975, n_29, n_28, n_1504, n_1490, n_1237, n_1236, n_1729, n_1728, n_1482;
  wire n_1336, n_1720, n_1330, n_939, n_1656, n_1439, n_1996, n_1997, n_1990, n_1991;
  wire n_1852, n_613, n_612, n_1721, n_1344, n_112, n_295, n_294, n_274, n_374;
  wire n_279, n_278, n_1576, n_1577, n_684, n_1548, n_206, n_1279, n_1278, n_1374;
  wire n_1273, n_1272, n_1925, n_1924, n_1888, n_1889, n_874, n_1077, n_1076, n_1880;
  wire n_50, n_51;
  assign n_0 = A[0];
  assign n_1 = A[0];
  assign n_2 = A[1];
  assign n_3 = A[1];
  assign n_4 = A[2];
  assign n_5 = A[2];
  assign n_6 = A[3];
  assign n_7 = A[3];
  assign n_8 = A[4];
  assign n_9 = A[4];
  assign n_10 = A[5];
  assign n_11 = A[5];
  assign n_12 = A[6];
  assign n_13 = A[6];
  assign n_14 = A[7];
  assign n_15 = A[7];
  assign n_16 = A[8];
  assign n_17 = A[8];
  assign n_18 = A[9];
  assign n_19 = A[9];
  assign n_20 = A[10];
  assign n_21 = A[10];
  assign n_22 = A[11];
  assign n_23 = A[11];
  assign n_24 = B[0];
  assign n_25 = B[0];
  assign n_26 = B[1];
  assign n_27 = B[1];
  assign n_28 = B[2];
  assign n_29 = B[2];
  assign n_30 = B[3];
  assign n_31 = B[3];
  assign n_32 = B[4];
  assign n_33 = B[4];
  assign n_34 = B[5];
  assign n_35 = B[5];
  assign n_36 = B[6];
  assign n_37 = B[6];
  assign n_38 = B[7];
  assign n_39 = B[7];
  assign n_40 = B[8];
  assign n_41 = B[8];
  assign n_42 = B[9];
  assign n_43 = B[9];
  assign n_44 = B[10];
  assign n_45 = B[10];
  assign n_46 = B[11];
  assign n_47 = B[11];
  assign n_50 = ~(n_38 & n_32 & n_42);
  assign n_51 = n_50;
  assign n_62 = ~(n_51 | n_32);
  assign n_63 = n_62;
  assign n_64 = ~(n_44 | n_28 | n_38);
  assign n_65 = n_64;
  assign n_66 = ~(n_65 & n_44 & n_22);
  assign n_70 = n_36 | n_66;
  assign n_71 = n_70;
  AOI21X1 tmp68(.Y(n_76), .A(n_2), .B(n_20), .C(n_71));
  assign n_77 = n_76;
  assign n_78 = ~(n_63 & n_62);
  assign n_104 = n_34 & n_28;
  assign n_105 = n_104;
  assign n_112 = n_105 & n_12;
  assign n_126 = n_22 & n_24;
  assign n_136 = ~(n_70 | n_70);
  assign n_137 = n_136;
  assign n_150 = ~n_137;
  assign n_184 = ~n_150;
  assign n_185 = n_184;
  assign n_206 = n_20 & n_26;
  assign n_214 = n_22 & n_26;
  assign n_228 = ~n_137;
  assign n_229 = n_228;
  assign n_230 = ~n_77;
  assign n_274 = ~n_230;
  assign n_278 = n_112 & n_32;
  assign n_279 = n_278;
  assign n_286 = ~(n_137 | n_150);
  assign n_287 = n_286;
  HAX1 tmp90(.YS(n_294), .YC(n_295), .A(n_126), .B(n_206));
  assign n_322 = n_295 & n_16;
  assign n_366 = n_18 & n_28;
  assign n_374 = n_20 & n_28;
  assign n_380 = n_22 & n_28;
  assign n_388 = ~(n_2 | n_78);
  assign n_416 = ~(n_2 | n_78);
  assign n_417 = n_416;
  assign n_428 = ~n_229;
  assign n_429 = n_428;
  FAX1 tmp100(.YS(n_452), .YC(n_453), .A(n_294), .B(n_366), .C(n_287));
  FAX1 tmp101(.YS(n_460), .YC(n_461), .A(n_214), .B(n_374), .C(n_295));
  assign n_518 = n_14 & n_30;
  assign n_526 = n_16 & n_30;
  assign n_532 = n_18 & n_30;
  assign n_540 = n_20 & n_30;
  assign n_548 = n_22 & n_30;
  assign n_604 = n_417 | n_518;
  assign n_605 = n_604;
  FAX1 tmp109(.YS(n_612), .YC(n_613), .A(n_452), .B(n_526), .C(n_279));
  FAX1 tmp110(.YS(n_620), .YC(n_621), .A(n_460), .B(n_532), .C(n_453));
  FAX1 tmp111(.YS(n_626), .YC(n_627), .A(n_380), .B(n_540), .C(n_461));
  assign n_684 = n_14 & n_32;
  assign n_692 = n_16 & n_32;
  assign n_700 = n_18 & n_32;
  assign n_706 = n_20 & n_32;
  assign n_714 = n_22 & n_32;
  assign n_764 = ~n_185;
  FAX1 tmp118(.YS(n_772), .YC(n_773), .A(n_612), .B(n_684), .C(n_605));
  FAX1 tmp119(.YS(n_778), .YC(n_779), .A(n_620), .B(n_692), .C(n_613));
  FAX1 tmp120(.YS(n_786), .YC(n_787), .A(n_626), .B(n_700), .C(n_621));
  FAX1 tmp121(.YS(n_794), .YC(n_795), .A(n_548), .B(n_706), .C(n_627));
  assign n_852 = n_14 & n_34;
  assign n_858 = n_16 & n_34;
  assign n_866 = n_18 & n_34;
  assign n_874 = n_20 & n_34;
  assign n_880 = n_22 & n_34;
  assign n_916 = ~(n_417 & n_28);
  assign n_917 = n_916;
  assign n_924 = ~(n_764 & n_274);
  assign n_925 = n_924;
  FAX1 tmp131(.YS(n_938), .YC(n_939), .A(n_778), .B(n_852), .C(n_773));
  FAX1 tmp132(.YS(n_946), .YC(n_947), .A(n_786), .B(n_858), .C(n_779));
  FAX1 tmp133(.YS(n_952), .YC(n_953), .A(n_794), .B(n_866), .C(n_787));
  FAX1 tmp134(.YS(n_960), .YC(n_961), .A(n_714), .B(n_874), .C(n_795));
  assign n_1004 = n_10 & n_36;
  assign n_1010 = n_12 & n_36;
  assign n_1018 = n_14 & n_36;
  assign n_1026 = n_16 & n_36;
  assign n_1032 = n_18 & n_36;
  assign n_1040 = n_20 & n_36;
  assign n_1048 = n_22 & n_36;
  assign n_1076 = ~n_137;
  assign n_1077 = n_1076;
  FAX1 tmp144(.YS(n_1084), .YC(n_1085), .A(n_924), .B(n_1010), .C(n_917));
  FAX1 tmp145(.YS(n_1090), .YC(n_1091), .A(n_63), .B(n_1004), .C(n_925));
  HAX1 tmp146(.YS(n_1098), .YC(n_1099), .A(n_938), .B(n_1010));
  FAX1 tmp147(.YS(n_1104), .YC(n_1105), .A(n_946), .B(n_1018), .C(n_939));
  FAX1 tmp148(.YS(n_1112), .YC(n_1113), .A(n_952), .B(n_1026), .C(n_947));
  FAX1 tmp149(.YS(n_1120), .YC(n_1121), .A(n_960), .B(n_1032), .C(n_953));
  FAX1 tmp150(.YS(n_1126), .YC(n_1127), .A(n_880), .B(n_1040), .C(n_961));
  assign n_1148 = n_4 & n_38;
  assign n_1162 = n_8 & n_38;
  assign n_1170 = n_10 & n_38;
  assign n_1178 = n_12 & n_38;
  assign n_1184 = n_14 & n_38;
  assign n_1192 = n_16 & n_38;
  assign n_1200 = n_18 & n_38;
  assign n_1206 = n_20 & n_38;
  assign n_1214 = n_22 & n_38;
  HAX1 tmp160(.YS(n_1236), .YC(n_1237), .A(n_1076), .B(n_1148));
  FAX1 tmp161(.YS(n_1242), .YC(n_1243), .A(n_1084), .B(n_150), .C(n_1077));
  FAX1 tmp162(.YS(n_1250), .YC(n_1251), .A(n_1090), .B(n_1162), .C(n_1085));
  FAX1 tmp163(.YS(n_1258), .YC(n_1259), .A(n_1098), .B(n_1170), .C(n_1091));
  FAX1 tmp164(.YS(n_1264), .YC(n_1265), .A(n_1104), .B(n_1178), .C(n_1099));
  FAX1 tmp165(.YS(n_1272), .YC(n_1273), .A(n_1112), .B(n_1184), .C(n_1105));
  FAX1 tmp166(.YS(n_1278), .YC(n_1279), .A(n_1120), .B(n_1192), .C(n_1113));
  FAX1 tmp167(.YS(n_1286), .YC(n_1287), .A(n_1126), .B(n_1200), .C(n_1121));
  FAX1 tmp168(.YS(n_1294), .YC(n_1295), .A(n_1048), .B(n_1206), .C(n_1127));
  assign n_1308 = n_2 & n_40;
  assign n_1316 = n_4 & n_40;
  assign n_1322 = n_6 & n_40;
  assign n_1330 = n_8 & n_40;
  assign n_1336 = n_10 & n_40;
  assign n_1344 = n_12 & n_40;
  assign n_1352 = n_14 & n_40;
  assign n_1358 = n_16 & n_40;
  assign n_1366 = n_18 & n_40;
  assign n_1374 = n_20 & n_40;
  assign n_1380 = n_22 & n_40;
  assign n_1394 = n_429 | n_1308;
  assign n_1395 = n_1394;
  FAX1 tmp182(.YS(n_1402), .YC(n_1403), .A(n_1242), .B(n_1316), .C(n_1237));
  FAX1 tmp183(.YS(n_1410), .YC(n_1411), .A(n_1250), .B(n_1322), .C(n_1243));
  FAX1 tmp184(.YS(n_1416), .YC(n_1417), .A(n_1258), .B(n_1330), .C(n_1251));
  FAX1 tmp185(.YS(n_1424), .YC(n_1425), .A(n_1264), .B(n_1336), .C(n_1259));
  FAX1 tmp186(.YS(n_1432), .YC(n_1433), .A(n_1272), .B(n_1344), .C(n_1265));
  FAX1 tmp187(.YS(n_1438), .YC(n_1439), .A(n_1278), .B(n_1352), .C(n_1273));
  FAX1 tmp188(.YS(n_1446), .YC(n_1447), .A(n_1286), .B(n_1358), .C(n_1279));
  FAX1 tmp189(.YS(n_1452), .YC(n_1453), .A(n_1294), .B(n_1366), .C(n_1287));
  FAX1 tmp190(.YS(n_1460), .YC(n_1461), .A(n_1214), .B(n_1374), .C(n_1295));
  assign n_1468 = n_0 & n_42;
  assign n_1482 = n_4 & n_42;
  assign n_1490 = n_6 & n_42;
  assign n_1496 = n_8 & n_42;
  assign n_1504 = n_10 & n_42;
  assign n_1510 = n_12 & n_42;
  assign n_1518 = n_14 & n_42;
  assign n_1526 = n_16 & n_42;
  assign n_1532 = n_18 & n_42;
  assign n_1540 = n_20 & n_42;
  assign n_1548 = n_22 & n_42;
  HAX1 tmp202(.YS(n_1554), .YC(n_1555), .A(n_6), .B(n_1468));
  FAX1 tmp203(.YS(n_1562), .YC(n_1563), .A(n_1402), .B(n_322), .C(n_1395));
  FAX1 tmp204(.YS(n_1568), .YC(n_1569), .A(n_1410), .B(n_1482), .C(n_1403));
  FAX1 tmp205(.YS(n_1576), .YC(n_1577), .A(n_1416), .B(n_1490), .C(n_1411));
  FAX1 tmp206(.YS(n_1584), .YC(n_1585), .A(n_1424), .B(n_1496), .C(n_1417));
  FAX1 tmp207(.YS(n_1590), .YC(n_1591), .A(n_1432), .B(n_1504), .C(n_1425));
  FAX1 tmp208(.YS(n_1598), .YC(n_1599), .A(n_1438), .B(n_1510), .C(n_1433));
  FAX1 tmp209(.YS(n_1604), .YC(n_1605), .A(n_1446), .B(n_1518), .C(n_1439));
  FAX1 tmp210(.YS(n_1612), .YC(n_1613), .A(n_1452), .B(n_1526), .C(n_1447));
  FAX1 tmp211(.YS(n_1620), .YC(n_1621), .A(n_1460), .B(n_1532), .C(n_1453));
  FAX1 tmp212(.YS(n_1626), .YC(n_1627), .A(n_1380), .B(n_1540), .C(n_1461));
  assign n_1634 = n_1555 & n_44;
  assign n_1642 = n_2 & n_44;
  assign n_1648 = n_4 & n_44;
  assign n_1656 = n_6 & n_44;
  assign n_1662 = n_8 & n_44;
  assign n_1670 = n_10 & n_44;
  assign n_1678 = n_12 & n_44;
  assign n_1684 = n_14 & n_44;
  assign n_1692 = n_16 & n_44;
  assign n_1700 = n_18 & n_44;
  assign n_1706 = n_20 & n_44;
  assign n_1714 = n_22 & n_44;
  FAX1 tmp225(.YS(n_1720), .YC(n_1721), .A(n_1562), .B(n_1634), .C(n_1555));
  FAX1 tmp226(.YS(n_1728), .YC(n_1729), .A(n_1568), .B(n_1642), .C(n_1563));
  FAX1 tmp227(.YS(n_1736), .YC(n_1737), .A(n_1576), .B(n_1648), .C(n_1569));
  FAX1 tmp228(.YS(n_1742), .YC(n_1743), .A(n_1584), .B(n_1656), .C(n_1577));
  FAX1 tmp229(.YS(n_1750), .YC(n_1751), .A(n_1590), .B(n_1662), .C(n_1585));
  FAX1 tmp230(.YS(n_1758), .YC(n_1759), .A(n_1598), .B(n_1670), .C(n_1591));
  FAX1 tmp231(.YS(n_1764), .YC(n_1765), .A(n_1604), .B(n_1678), .C(n_1599));
  FAX1 tmp232(.YS(n_1772), .YC(n_1773), .A(n_1612), .B(n_1684), .C(n_1605));
  FAX1 tmp233(.YS(n_1778), .YC(n_1779), .A(n_1620), .B(n_1692), .C(n_1613));
  FAX1 tmp234(.YS(n_1786), .YC(n_1787), .A(n_1626), .B(n_1700), .C(n_1621));
  FAX1 tmp235(.YS(n_1794), .YC(n_1795), .A(n_1548), .B(n_1706), .C(n_1627));
  assign n_1800 = n_0 & n_46;
  assign n_1808 = n_2 & n_46;
  assign n_1816 = n_4 & n_46;
  assign n_1822 = n_6 & n_46;
  assign n_1830 = n_8 & n_46;
  assign n_1836 = n_10 & n_46;
  assign n_1844 = n_12 & n_46;
  assign n_1852 = n_14 & n_46;
  assign n_1858 = n_16 & n_46;
  assign n_1866 = n_18 & n_46;
  assign n_1874 = n_20 & n_46;
  assign n_1880 = n_22 & n_46;
  FAX1 tmp248(.YS(n_1888), .YC(n_1889), .A(n_1728), .B(n_1800), .C(n_1721));
  FAX1 tmp249(.YS(n_1894), .YC(n_1895), .A(n_1736), .B(n_1808), .C(n_1729));
  FAX1 tmp250(.YS(n_1902), .YC(n_1903), .A(n_1742), .B(n_1816), .C(n_1737));
  FAX1 tmp251(.YS(n_1910), .YC(n_1911), .A(n_1750), .B(n_1822), .C(n_1743));
  FAX1 tmp252(.YS(n_1916), .YC(n_1917), .A(n_1758), .B(n_1830), .C(n_1751));
  FAX1 tmp253(.YS(n_1924), .YC(n_1925), .A(n_1764), .B(n_1836), .C(n_1759));
  FAX1 tmp254(.YS(n_1932), .YC(n_1933), .A(n_1772), .B(n_1844), .C(n_1765));
  FAX1 tmp255(.YS(n_1938), .YC(n_1939), .A(n_1778), .B(n_1852), .C(n_1773));
  FAX1 tmp256(.YS(n_1946), .YC(n_1947), .A(n_1786), .B(n_1858), .C(n_1779));
  FAX1 tmp257(.YS(n_1952), .YC(n_1953), .A(n_1794), .B(n_1866), .C(n_1787));
  FAX1 tmp258(.YS(n_1960), .YC(n_1961), .A(n_1714), .B(n_1874), .C(n_1795));
  HAX1 tmp259(.YS(n_1968), .YC(n_1969), .A(n_1894), .B(n_1889));
  FAX1 tmp260(.YS(n_1974), .YC(n_1975), .A(n_1902), .B(n_1895), .C(n_1969));
  FAX1 tmp261(.YS(n_1982), .YC(n_1983), .A(n_1910), .B(n_1903), .C(n_1975));
  FAX1 tmp262(.YS(n_1990), .YC(n_1991), .A(n_1916), .B(n_1911), .C(n_1983));
  FAX1 tmp263(.YS(n_1996), .YC(n_1997), .A(n_1924), .B(n_1917), .C(n_1991));
  FAX1 tmp264(.YS(n_2004), .YC(n_2005), .A(n_1932), .B(n_1925), .C(n_1997));
  FAX1 tmp265(.YS(n_2010), .YC(n_2011), .A(n_1938), .B(n_1933), .C(n_2005));
  FAX1 tmp266(.YS(n_2018), .YC(n_2019), .A(n_1946), .B(n_1939), .C(n_2011));
  FAX1 tmp267(.YS(n_2026), .YC(n_2027), .A(n_1952), .B(n_1947), .C(n_2019));
  FAX1 tmp268(.YS(n_2032), .YC(n_2033), .A(n_1960), .B(n_1953), .C(n_2027));
  FAX1 tmp269(.YS(n_2040), .YC(n_2041), .A(n_1880), .B(n_1961), .C(n_2033));
  assign O[0] = n_953;
  assign O[1] = n_78;
  assign O[2] = n_388;
  assign O[3] = n_0;
  assign O[4] = n_429;
  assign O[5] = n_66;
  assign O[6] = n_287;
  assign O[7] = n_916;
  assign O[8] = n_34;
  assign O[9] = n_1554;
  assign O[10] = n_1720;
  assign O[11] = n_1888;
  assign O[12] = n_1968;
  assign O[13] = n_1974;
  assign O[14] = n_1982;
  assign O[15] = n_1990;
  assign O[16] = n_1996;
  assign O[17] = n_2004;
  assign O[18] = n_2010;
  assign O[19] = n_2018;
  assign O[20] = n_2026;
  assign O[21] = n_2032;
  assign O[22] = n_2040;
  assign O[23] = n_2041;
endmodule


// internal reference: cgp-compare17.12.mul12u_pwr_0_680_wce_00_0493

