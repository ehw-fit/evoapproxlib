/***
* This code is a part of ApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under a XXXX public license.
* When used, please cite the following article: tbd 
* This file is pareto optimal sub-set in the pwr and wce parameters
***/

module mul12u_pwr_0_028_wce_09_7620(A, B, O);
  input [11:0] A, B;
  output [23:0] O;
  wire n_1274, n_1049, n_42, n_1287, n_1285, n_1283, n_1281, n_1289, n_1051, n_1180;
  wire n_1420, n_1182, n_1512, n_1510, n_1516, n_1514, n_1518, n_1027, n_1024, n_23;
  wire n_22, n_21, n_20, n_920, n_25, n_29, n_1500, n_1502, n_129, n_1504;
  wire n_1506, n_1508, n_650, n_1408, n_1400, n_0, n_1402, n_1404, n_1406, n_1484;
  wire n_422, n_18, n_19, n_16, n_17, n_14, n_15, n_12, n_13, n_10;
  wire n_11, n_1158, n_1498, n_1152, n_1150, n_1494, n_1156, n_1490, n_81, n_1522;
  wire n_1520, n_1012, n_1311, n_1313, n_1393, n_1395, n_71, n_1416, n_1414, n_213;
  wire n_1412, n_1410, n_1418, n_1307, n_566, n_1178, n_1309, n_8, n_9, n_4;
  wire n_5, n_6, n_7, n_1277, n_1, n_2, n_3;
  assign n_0 = A[0];
  assign n_1 = A[1];
  assign n_2 = A[2];
  assign n_3 = A[3];
  assign n_4 = A[4];
  assign n_5 = A[5];
  assign n_6 = A[6];
  assign n_7 = A[7];
  assign n_8 = A[8];
  assign n_9 = A[9];
  assign n_10 = A[10];
  assign n_11 = A[11];
  assign n_12 = B[0];
  assign n_13 = B[1];
  assign n_14 = B[2];
  assign n_15 = B[3];
  assign n_16 = B[4];
  assign n_17 = B[5];
  assign n_18 = B[6];
  assign n_19 = B[7];
  assign n_20 = B[8];
  assign n_21 = B[9];
  assign n_22 = B[10];
  assign n_23 = B[11];
  assign n_25 = ~(n_18 | n_17);
  assign n_29 = n_25 & n_18;
  assign n_42 = ~n_29;
  assign n_71 = n_42;
  assign n_81 = n_23 & n_21;
  assign n_129 = ~(n_29 | n_71);
  assign n_213 = n_19 & n_29;
  assign n_422 = ~n_29;
  assign n_566 = ~n_129;
  assign n_650 = ~n_71;
  assign n_920 = n_11 & n_20;
  assign n_1012 = n_29 & n_422;
  assign n_1024 = n_81 & n_10;
  assign n_1027 = n_1012 | n_1024;
  assign n_1049 = n_10 & n_21;
  assign n_1051 = n_11 & n_21;
  assign n_1150 = n_920 ^ n_650;
  assign n_1152 = n_920 & n_1049;
  assign n_1156 = n_1150 | n_1027;
  assign n_1158 = n_1152 | n_1012;
  assign n_1178 = n_9 & n_22;
  assign n_1180 = n_10 & n_22;
  assign n_1182 = n_11 & n_22;
  assign n_1274 = n_1156 & n_1178;
  assign n_1277 = ~(n_650 | n_422);
  assign n_1281 = n_1051 ^ n_1180;
  assign n_1283 = n_1051 & n_1180;
  assign n_1285 = n_20 & n_1158;
  assign n_1287 = n_1281 ^ n_1158;
  assign n_1289 = n_1283 | n_1285;
  assign n_1307 = n_8 & n_23;
  assign n_1309 = n_9 & n_23;
  assign n_1311 = n_10 & n_23;
  assign n_1313 = n_11 & n_23;
  assign n_1393 = n_129 ^ n_1307;
  assign n_1395 = ~n_1277;
  assign n_1400 = n_213;
  assign n_1402 = n_1287 ^ n_1309;
  assign n_1404 = n_1287 & n_1309;
  assign n_1406 = n_1402 & n_1274;
  assign n_1408 = n_1402 ^ n_1274;
  assign n_1410 = n_1404 | n_1406;
  assign n_1412 = n_1182 ^ n_1311;
  assign n_1414 = n_1182 & n_1311;
  assign n_1416 = n_1412 & n_1289;
  assign n_1418 = n_1412 ^ n_1289;
  assign n_1420 = n_1414 | n_1416;
  assign n_1484 = n_1393 ^ n_422;
  assign n_1490 = ~n_1484;
  assign n_1494 = n_1408 ^ n_1400;
  assign n_1498 = n_1494 & n_566;
  assign n_1500 = n_1494 ^ n_566;
  assign n_1502 = n_129 | n_1498;
  assign n_1504 = n_1418 ^ n_1410;
  assign n_1506 = n_1418 & n_1410;
  assign n_1508 = n_1504 & n_1494;
  assign n_1510 = n_1504 ^ n_1502;
  assign n_1512 = n_1506 | n_1508;
  assign n_1514 = n_1313 ^ n_1420;
  assign n_1516 = n_1313 & n_1420;
  assign n_1518 = n_1514 & n_1512;
  assign n_1520 = n_1514 ^ n_1512;
  assign n_1522 = n_1516 | n_1518;
  assign O[0] = n_13;
  assign O[1] = n_6;
  assign O[2] = n_1395;
  assign O[3] = n_1012;
  assign O[4] = n_17;
  assign O[5] = n_18;
  assign O[6] = n_7;
  assign O[7] = n_1400;
  assign O[8] = n_129;
  assign O[9] = n_2;
  assign O[10] = n_19;
  assign O[11] = n_16;
  assign O[12] = n_1;
  assign O[13] = n_422;
  assign O[14] = n_23;
  assign O[15] = n_4;
  assign O[16] = n_21;
  assign O[17] = n_6;
  assign O[18] = n_7;
  assign O[19] = n_1490;
  assign O[20] = n_1500;
  assign O[21] = n_1510;
  assign O[22] = n_1520;
  assign O[23] = n_1522;
endmodule


// internal reference: cgp-compare17.12.mul12u_pwr_0_028_wce_09_7620

