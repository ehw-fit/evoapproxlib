/***
* This code is a part of ApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under a XXXX public license.
* When used, please cite the following article: tbd 
* This file is pareto optimal sub-set in the pdk45_pwr and mae% parameters
***/

// ../../../cgp.nn/res/11b_160129\wtm_rca\e15.0\run.00376.txt
module mul11u_pwr_0_084_mae_03_3411(A, B, O);
  input [10:0] A, B;
  output [21:0] O;
  wire [10:0] A, B;
  wire [21:0] O;
  wire sig_65, sig_75, sig_99, sig_105, sig_108, sig_109;
  wire sig_115, sig_118, sig_119, sig_120, sig_123, sig_128;
  wire sig_129, sig_130, sig_131, sig_133, sig_139, sig_140;
  wire sig_142, sig_198, sig_234, sig_256, sig_264, sig_267;
  wire sig_268, sig_271, sig_279, sig_282, sig_283, sig_284;
  wire sig_285, sig_286, sig_287, sig_288, sig_343, sig_357;
  wire sig_358, sig_360, sig_371, sig_386, sig_387, sig_388;
  wire sig_389, sig_390, sig_391, sig_406, sig_409, sig_452;
  wire sig_478, sig_481, sig_482, sig_483, sig_484, sig_485;
  wire sig_486, sig_487, sig_488, sig_489, sig_490, sig_491;
  wire sig_492, sig_493, sig_494, sig_495, sig_496, sig_504;
  wire sig_505, sig_547, sig_549, sig_550, sig_552, sig_553;
  wire sig_554, sig_555, sig_556, sig_598, sig_601, sig_602;
  wire sig_603, sig_605, sig_606, sig_607, sig_608, sig_609;
  wire sig_610, sig_611, sig_612, sig_613, sig_614, sig_615;
  wire sig_616, sig_617, sig_671, sig_672, sig_673, sig_675;
  wire sig_676, sig_677, sig_678, sig_680, sig_681, sig_682;
  wire sig_683, sig_685, sig_686, sig_687, sig_688, sig_690;
  assign O[12] = A[10] & B[1];
  assign O[16] = A[1] & B[3];
  assign sig_65 = A[4] & B[1];
  assign sig_75 = A[6] & B[4];
  assign O[15] = A[4] & B[6];
  assign sig_99 = A[3] & B[7];
  assign sig_105 = B[6] & B[7];
  assign sig_108 = A[9] & B[7];
  assign sig_109 = A[10] & B[7];
  assign sig_115 = B[0] ^ B[9];
  assign sig_118 = A[4] & B[2];
  assign sig_119 = A[9] & B[8];
  assign sig_120 = A[10] & B[8];
  assign sig_123 = A[2] & B[9];
  assign sig_128 = A[7] & A[9];
  assign sig_129 = A[8] & B[9];
  assign sig_130 = A[9] & B[9];
  assign sig_131 = A[10] & B[9];
  assign sig_133 = A[1] & B[10];
  assign O[4] = A[2] & B[10];
  assign sig_139 = A[7] & B[10];
  assign sig_140 = A[8] & B[10];
  assign O[2] = A[9] & B[10];
  assign sig_142 = A[10] & B[10];
  assign O[13] = O[16] & A[1];
  assign sig_198 = B[10] | B[10];
  assign O[5] = A[2] & B[10];
  assign sig_234 = sig_65 ^ sig_75;
  assign O[11] = sig_234;
  assign O[9] = B[9] & sig_99;
  assign sig_256 = B[1];
  assign sig_264 = A[2];
  assign sig_267 = sig_264;
  assign sig_268 = B[4] ^ sig_105;
  assign sig_271 = sig_268 ^ sig_115;
  assign sig_279 = !(B[9] | B[10]);
  assign sig_282 = sig_279;
  assign sig_283 = O[15];
  assign sig_284 = O[15] ^ sig_108;
  assign sig_285 = B[9] & A[7];
  assign sig_286 = sig_283 ^ sig_118;
  assign sig_287 = sig_284 | sig_285;
  assign sig_288 = sig_109 & sig_119;
  assign O[0] = sig_109 ^ sig_119;
  assign O[8] = B[4] & A[3];
  assign sig_343 = sig_198 & B[1];
  assign sig_357 = A[10] & sig_256;
  assign sig_358 = A[3] & B[7];
  assign sig_360 = sig_357 | sig_358;
  assign sig_371 = B[2] ^ sig_271;
  assign O[10] = sig_371 & sig_267;
  assign sig_386 = sig_286 & sig_282;
  assign sig_387 = sig_286 ^ B[6];
  assign sig_388 = O[0] & sig_287;
  assign sig_389 = O[0] ^ sig_287;
  assign sig_390 = sig_120 & sig_288;
  assign sig_391 = sig_120 ^ sig_288;
  assign sig_406 = B[7] & A[7];
  assign sig_409 = sig_406;
  assign sig_452 = sig_360 ^ sig_123;
  assign O[1] = sig_452 ^ sig_133;
  assign sig_478 = B[2] & sig_128;
  assign sig_481 = sig_478;
  assign sig_482 = sig_386 ^ sig_129;
  assign sig_483 = sig_386 & sig_129;
  assign sig_484 = sig_482 & sig_139;
  assign sig_485 = sig_482 ^ sig_139;
  assign sig_486 = sig_483 | sig_484;
  assign sig_487 = sig_388 ^ sig_130;
  assign sig_488 = sig_388 & sig_130;
  assign sig_489 = sig_487 & sig_140;
  assign sig_490 = sig_487 ^ sig_140;
  assign sig_491 = sig_488 ^ sig_489;
  assign sig_492 = sig_390 ^ sig_131;
  assign sig_493 = sig_390 & sig_131;
  assign sig_494 = sig_492 & O[2];
  assign sig_495 = sig_492 ^ O[2];
  assign sig_496 = sig_493 | sig_494;
  assign sig_504 = sig_409;
  assign sig_505 = A[2] & sig_343;
  assign O[3] = sig_504 | sig_505;
  assign sig_547 = B[5];
  assign sig_549 = sig_387 & A[4];
  assign sig_550 = B[10] & A[9];
  assign sig_552 = sig_549 | sig_550;
  assign sig_553 = sig_389 & sig_485;
  assign sig_554 = sig_389 ^ sig_485;
  assign sig_555 = sig_391 & sig_490;
  assign sig_556 = sig_391 ^ sig_490;
  assign O[7] = B[6] & A[2];
  assign sig_598 = A[7] & sig_547;
  assign sig_601 = sig_598;
  assign sig_602 = sig_554 ^ sig_552;
  assign sig_603 = B[8] & sig_552;
  assign sig_605 = sig_602 ^ sig_481;
  assign sig_606 = sig_603;
  assign sig_607 = sig_556 ^ sig_553;
  assign sig_608 = sig_556 & sig_553;
  assign sig_609 = sig_607 & sig_486;
  assign sig_610 = sig_607 ^ sig_486;
  assign sig_611 = sig_608 | sig_609;
  assign sig_612 = sig_495 ^ sig_555;
  assign sig_613 = sig_495 & sig_555;
  assign sig_614 = sig_612 & sig_491;
  assign sig_615 = sig_612 ^ sig_491;
  assign sig_616 = sig_613 | sig_614;
  assign sig_617 = sig_142 & sig_496;
  assign O[14] = sig_142 ^ sig_496;
  assign sig_671 = sig_605 ^ sig_601;
  assign sig_672 = sig_605 & sig_601;
  assign sig_673 = sig_671 & A[6];
  assign sig_675 = sig_672 & sig_673;
  assign sig_676 = sig_610 ^ sig_606;
  assign sig_677 = sig_610 & sig_606;
  assign sig_678 = A[1] & sig_675;
  assign O[18] = sig_676 ^ sig_675;
  assign sig_680 = sig_677 | sig_678;
  assign sig_681 = sig_615 ^ sig_611;
  assign sig_682 = sig_615 & sig_611;
  assign sig_683 = sig_681 & sig_680;
  assign O[19] = sig_681 ^ sig_680;
  assign sig_685 = sig_682 | sig_683;
  assign sig_686 = O[14] ^ sig_616;
  assign sig_687 = O[14] & sig_616;
  assign sig_688 = sig_686 & sig_685;
  assign O[20] = sig_686 ^ sig_685;
  assign sig_690 = sig_687 | sig_688;
  assign O[21] = sig_617 ^ sig_690;
  assign O[6] = O[1]; // default output
  assign O[17] = O[5]; // default output
endmodule


// internal reference: cgp-nn-iccad16.11.mul11u_pwr_0_084_mae_03_3411

