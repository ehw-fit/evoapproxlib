/***
* This code is a part of ApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under a XXXX public license.
* When used, please cite the following article: tbd 
* This file is pareto optimal sub-set in the pdk45_pwr and ep% parameters
***/

// ../../../cgp.nn/res/7b_160129\rcam\e00.5\run.00686.txt
module mul7u_pwr_0_208_ep_91(A, B, O);
  input [6:0] A, B;
  output [13:0] O;
  wire [6:0] A, B;
  wire [13:0] O;
  wire sig_19, sig_20, sig_25, sig_26, sig_27, sig_45;
  wire sig_46, sig_48, sig_49, sig_50, sig_51, sig_52;
  wire sig_53, sig_54, sig_55, sig_56, sig_61, sig_62;
  wire sig_63, sig_76, sig_79, sig_80, sig_81, sig_82;
  wire sig_83, sig_84, sig_85, sig_86, sig_87, sig_88;
  wire sig_89, sig_90, sig_91, sig_92, sig_93, sig_95;
  wire sig_98, sig_99, sig_100, sig_101, sig_102, sig_110;
  wire sig_111, sig_113, sig_114, sig_115, sig_116, sig_117;
  wire sig_118, sig_119, sig_120, sig_121, sig_122, sig_123;
  wire sig_124, sig_125, sig_126, sig_127, sig_128, sig_129;
  wire sig_130, sig_131, sig_132, sig_133, sig_136, sig_137;
  wire sig_138, sig_139, sig_140, sig_141, sig_144, sig_145;
  wire sig_147, sig_148, sig_149, sig_150, sig_151, sig_152;
  wire sig_153, sig_154, sig_156, sig_157, sig_158, sig_159;
  wire sig_160, sig_161, sig_162, sig_163, sig_164, sig_165;
  wire sig_166, sig_167, sig_168, sig_169, sig_170, sig_171;
  wire sig_172, sig_173, sig_174, sig_175, sig_176, sig_177;
  wire sig_178, sig_179, sig_180, sig_182, sig_183, sig_184;
  wire sig_185, sig_186, sig_187, sig_188, sig_189, sig_190;
  wire sig_191, sig_192, sig_193, sig_194, sig_195, sig_196;
  wire sig_197, sig_198, sig_199, sig_200, sig_201, sig_202;
  wire sig_203, sig_204, sig_205, sig_206, sig_207, sig_208;
  wire sig_209, sig_210, sig_211, sig_212, sig_214, sig_215;
  wire sig_216, sig_217, sig_218, sig_219, sig_221, sig_222;
  wire sig_223, sig_224, sig_226, sig_227, sig_228, sig_229;
  wire sig_231, sig_232, sig_233, sig_236, sig_237, sig_238;
  wire sig_239, sig_241, sig_242, sig_243, sig_244, sig_246;
  wire sig_247, sig_248, sig_249;
  assign sig_19 = A[5] & B[0];
  assign sig_20 = A[6] & B[0];
  assign sig_25 = A[4] & B[1];
  assign sig_26 = A[5] & B[1];
  assign sig_27 = A[6] & B[1];
  assign sig_45 = sig_19 ^ sig_25;
  assign sig_46 = A[5] & A[4];
  assign sig_48 = sig_45;
  assign sig_49 = sig_46 & B[1];
  assign sig_50 = sig_20 ^ sig_26;
  assign sig_51 = sig_20 & sig_26;
  assign sig_52 = B[0] & sig_49;
  assign sig_53 = sig_50 | sig_49;
  assign sig_54 = sig_51 | sig_52;
  assign sig_55 = sig_54 ^ sig_27;
  assign sig_56 = sig_54 & A[6];
  assign sig_61 = A[4] & B[2];
  assign sig_62 = A[5] & B[2];
  assign sig_63 = A[6] & B[2];
  assign sig_76 = sig_48;
  assign sig_79 = sig_76;
  assign sig_80 = B[2] & A[3];
  assign sig_81 = sig_53 ^ sig_61;
  assign sig_82 = sig_53 & sig_61;
  assign sig_83 = sig_81 & sig_80;
  assign sig_84 = sig_81 ^ sig_80;
  assign sig_85 = sig_82 ^ sig_83;
  assign sig_86 = sig_55 ^ sig_62;
  assign sig_87 = sig_55 & sig_62;
  assign sig_88 = sig_86 & sig_85;
  assign sig_89 = sig_86 ^ sig_85;
  assign sig_90 = sig_87 ^ sig_88;
  assign sig_91 = sig_56 ^ sig_63;
  assign sig_92 = sig_56 & B[2];
  assign sig_93 = A[6] & sig_90;
  assign O[0] = sig_91 ^ sig_90;
  assign sig_95 = sig_92 | sig_93;
  assign sig_98 = A[2] & B[3];
  assign sig_99 = A[3] & B[3];
  assign sig_100 = A[4] & B[3];
  assign sig_101 = A[5] & B[3];
  assign sig_102 = A[6] & B[3];
  assign sig_110 = sig_79 | sig_98;
  assign sig_111 = sig_79 & A[2];
  assign sig_113 = sig_110;
  assign sig_114 = sig_111 & B[3];
  assign sig_115 = sig_84 ^ sig_99;
  assign sig_116 = sig_84 & sig_99;
  assign sig_117 = sig_115 & sig_114;
  assign sig_118 = sig_115 ^ sig_114;
  assign sig_119 = sig_116 | sig_117;
  assign sig_120 = sig_89 ^ sig_100;
  assign sig_121 = sig_89 & sig_100;
  assign sig_122 = sig_120 & sig_119;
  assign sig_123 = sig_120 ^ sig_119;
  assign sig_124 = sig_121 | sig_122;
  assign sig_125 = O[0] ^ sig_101;
  assign sig_126 = O[0] & sig_101;
  assign sig_127 = sig_125 & sig_124;
  assign sig_128 = sig_125 ^ sig_124;
  assign sig_129 = sig_126 ^ sig_127;
  assign sig_130 = sig_95 ^ sig_102;
  assign sig_131 = sig_95 & B[3];
  assign sig_132 = A[6] & sig_129;
  assign sig_133 = sig_130 ^ sig_129;
  assign O[3] = sig_131 | sig_132;
  assign sig_136 = A[1] & B[4];
  assign sig_137 = A[2] & B[4];
  assign sig_138 = A[3] & B[4];
  assign sig_139 = A[4] & B[4];
  assign sig_140 = A[5] & B[4];
  assign sig_141 = A[6] & B[4];
  assign sig_144 = sig_113 | sig_136;
  assign sig_145 = sig_113 & A[1];
  assign sig_147 = sig_144;
  assign sig_148 = sig_145 & B[4];
  assign sig_149 = sig_118 ^ sig_137;
  assign sig_150 = sig_118 & sig_137;
  assign sig_151 = sig_149 & sig_148;
  assign sig_152 = sig_149 ^ sig_148;
  assign sig_153 = sig_150 ^ sig_151;
  assign sig_154 = sig_123 ^ sig_138;
  assign O[1] = sig_123 & sig_138;
  assign sig_156 = sig_154 & sig_153;
  assign sig_157 = sig_154 ^ sig_153;
  assign sig_158 = O[1] | sig_156;
  assign sig_159 = sig_128 ^ sig_139;
  assign sig_160 = sig_128 & sig_139;
  assign sig_161 = sig_159 & sig_158;
  assign sig_162 = sig_159 ^ sig_158;
  assign sig_163 = sig_160 ^ sig_161;
  assign sig_164 = sig_133 ^ sig_140;
  assign sig_165 = sig_133 & sig_140;
  assign sig_166 = sig_164 & sig_163;
  assign sig_167 = sig_164 ^ sig_163;
  assign sig_168 = sig_165 ^ sig_166;
  assign sig_169 = O[3] ^ sig_141;
  assign sig_170 = O[3] & B[4];
  assign sig_171 = A[6] & sig_168;
  assign sig_172 = sig_169 ^ sig_168;
  assign sig_173 = sig_170 | sig_171;
  assign sig_174 = A[0] & B[5];
  assign sig_175 = A[1] & B[5];
  assign sig_176 = A[2] & B[5];
  assign sig_177 = A[3] & B[5];
  assign sig_178 = A[4] & B[5];
  assign sig_179 = A[5] & B[5];
  assign sig_180 = A[6] & B[5];
  assign O[5] = sig_147 | sig_174;
  assign sig_182 = sig_147 & sig_174;
  assign sig_183 = sig_152 ^ sig_175;
  assign sig_184 = sig_152 & sig_175;
  assign sig_185 = sig_183 & sig_182;
  assign sig_186 = sig_183 ^ sig_182;
  assign sig_187 = sig_184 | sig_185;
  assign sig_188 = sig_157 ^ sig_176;
  assign sig_189 = sig_157 & sig_176;
  assign sig_190 = sig_188 & sig_187;
  assign sig_191 = sig_188 ^ sig_187;
  assign sig_192 = sig_189 | sig_190;
  assign sig_193 = sig_162 ^ sig_177;
  assign sig_194 = sig_162 & sig_177;
  assign sig_195 = sig_193 & sig_192;
  assign sig_196 = sig_193 ^ sig_192;
  assign sig_197 = sig_194 | sig_195;
  assign sig_198 = sig_167 ^ sig_178;
  assign sig_199 = sig_167 & sig_178;
  assign sig_200 = sig_198 & sig_197;
  assign sig_201 = sig_198 ^ sig_197;
  assign sig_202 = sig_199 | sig_200;
  assign sig_203 = sig_172 ^ sig_179;
  assign sig_204 = sig_172 & sig_179;
  assign sig_205 = sig_203 & sig_202;
  assign sig_206 = sig_203 ^ sig_202;
  assign sig_207 = sig_204 | sig_205;
  assign sig_208 = sig_173 ^ sig_180;
  assign sig_209 = sig_173 & B[5];
  assign sig_210 = A[6] & sig_207;
  assign sig_211 = sig_208 ^ sig_207;
  assign sig_212 = sig_209 | sig_210;
  assign O[4] = A[0] & B[6];
  assign sig_214 = A[1] & B[6];
  assign sig_215 = A[2] & B[6];
  assign sig_216 = A[3] & B[6];
  assign sig_217 = A[4] & B[6];
  assign sig_218 = A[5] & B[6];
  assign sig_219 = A[6] & B[6];
  assign O[6] = sig_186 ^ O[4];
  assign sig_221 = sig_186 & O[4];
  assign sig_222 = sig_191 ^ sig_214;
  assign sig_223 = sig_191 & sig_214;
  assign sig_224 = sig_222 & sig_221;
  assign O[7] = sig_222 ^ sig_221;
  assign sig_226 = sig_223 | sig_224;
  assign sig_227 = sig_196 ^ sig_215;
  assign sig_228 = sig_196 & sig_215;
  assign sig_229 = sig_227 & sig_226;
  assign O[8] = sig_227 ^ sig_226;
  assign sig_231 = sig_228 ^ sig_229;
  assign sig_232 = sig_201 ^ sig_216;
  assign sig_233 = sig_201 & sig_216;
  assign O[2] = sig_232 & sig_231;
  assign O[9] = sig_232 ^ sig_231;
  assign sig_236 = sig_233 | O[2];
  assign sig_237 = sig_206 ^ sig_217;
  assign sig_238 = sig_206 & sig_217;
  assign sig_239 = sig_237 & sig_236;
  assign O[10] = sig_237 ^ sig_236;
  assign sig_241 = sig_238 | sig_239;
  assign sig_242 = sig_211 ^ sig_218;
  assign sig_243 = sig_211 & sig_218;
  assign sig_244 = sig_242 & sig_241;
  assign O[11] = sig_242 ^ sig_241;
  assign sig_246 = sig_243 | sig_244;
  assign sig_247 = sig_212 ^ sig_219;
  assign sig_248 = sig_212 & B[6];
  assign sig_249 = A[6] & sig_246;
  assign O[12] = sig_247 ^ sig_246;
  assign O[13] = sig_248 | sig_249;
endmodule


// internal reference: cgp-nn-iccad16.07.mul7u_pwr_0_208_ep_91

