/***
    * This code is a part of ApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under a XXXX public license.
    * When used, please cite the following article: tbd 
    * This file is pareto optimal sub-set in the pwr and mae parameters
    ***/
    
module mul12u_pwr_0_427_mae_00_0729(A, B, O);
  input [11:0] A, B;
  output [23:0] O;
  wire n_947, n_946, n_548, n_1947, n_1366, n_704, n_707, n_706, n_1192, n_700;
  wire n_45, n_44, n_47, n_46, n_41, n_40, n_43, n_42, n_1040, n_1759;
  wire n_866, n_1591, n_49, n_48, n_1200, n_1286, n_380, n_2018, n_2019, n_1874;
  wire n_1743, n_2010, n_2011, n_1742, n_778, n_779, n_1786, n_2027, n_1684, n_1446;
  wire n_1447, n_1295, n_952, n_540, n_1358, n_1621, n_1214, n_1294, n_1184, n_714;
  wire n_1425, n_1352, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37;
  wire n_38, n_39, n_1585, n_1584, n_392, n_393, n_1991, n_1751, n_1787, n_152;
  wire n_153, n_2005, n_787, n_156, n_157, n_1121, n_1510, n_786, n_1952, n_1453;
  wire n_1112, n_1518, n_1933, n_1113, n_1953, n_1026, n_1438, n_1120, n_1344, n_23;
  wire n_22, n_21, n_20, n_27, n_26, n_25, n_24, n_1974, n_29, n_28;
  wire n_1336, n_1590, n_1866, n_1613, n_1612, n_1598, n_1273, n_1692, n_1946, n_1504;
  wire n_1272, n_127, n_126, n_1032, n_1287, n_1982, n_1642, n_1822, n_932, n_933;
  wire n_18, n_19, n_16, n_17, n_14, n_15, n_12, n_13, n_10, n_11;
  wire n_1758, n_648, n_649, n_880, n_1844, n_136, n_137, n_2033, n_1532, n_2026;
  wire n_1714, n_626, n_627, n_620, n_621, n_1127, n_1656, n_1126, n_1439, n_1961;
  wire n_1491, n_1490, n_1996, n_1960, n_1916, n_1917, n_1910, n_1911, n_532, n_1997;
  wire n_1627, n_938, n_1048, n_1858, n_2032, n_939, n_1526, n_1054, n_1018, n_1548;
  wire n_1259, n_1258, n_1010, n_1540, n_1620, n_692, n_1662, n_1433, n_853, n_852;
  wire n_1099, n_1098, n_858, n_1902, n_2041, n_2040, n_1903, n_1852, n_215, n_214;
  wire n_1983, n_1706, n_1794, n_1795, n_1176, n_270, n_1264, n_1265, n_1678, n_1178;
  wire n_1626, n_1599, n_953, n_1772, n_1773, n_1452, n_961, n_960, n_1778, n_1670;
  wire n_1938, n_1939, n_2004, n_1750, n_1388, n_280, n_281, n_65, n_64, n_1206;
  wire n_1380, n_994, n_995, n_1460, n_1461, n_1830, n_1779, n_1432, n_1424, n_1837;
  wire n_1836, n_1279, n_1278, n_8, n_9, n_1374, n_4, n_5, n_6, n_7;
  wire n_0, n_1, n_2, n_3, n_1765, n_1764, n_1925, n_1924, n_874, n_1880;
  wire n_1604, n_1605, n_1105, n_1990, n_1104, n_794, n_54, n_795, n_1700, n_1932;
  wire n_761, n_760;
  assign n_0 = A[0];
  assign n_1 = A[0];
  assign n_2 = A[1];
  assign n_3 = A[1];
  assign n_4 = A[2];
  assign n_5 = A[2];
  assign n_6 = A[3];
  assign n_7 = A[3];
  assign n_8 = A[4];
  assign n_9 = A[4];
  assign n_10 = A[5];
  assign n_11 = A[5];
  assign n_12 = A[6];
  assign n_13 = A[6];
  assign n_14 = A[7];
  assign n_15 = A[7];
  assign n_16 = A[8];
  assign n_17 = A[8];
  assign n_18 = A[9];
  assign n_19 = A[9];
  assign n_20 = A[10];
  assign n_21 = A[10];
  assign n_22 = A[11];
  assign n_23 = A[11];
  assign n_24 = B[0];
  assign n_25 = B[0];
  assign n_26 = B[1];
  assign n_27 = B[1];
  assign n_28 = B[2];
  assign n_29 = B[2];
  assign n_30 = B[3];
  assign n_31 = B[3];
  assign n_32 = B[4];
  assign n_33 = B[4];
  assign n_34 = B[5];
  assign n_35 = B[5];
  assign n_36 = B[6];
  assign n_37 = B[6];
  assign n_38 = B[7];
  assign n_39 = B[7];
  assign n_40 = B[8];
  assign n_41 = B[8];
  assign n_42 = B[9];
  assign n_43 = B[9];
  assign n_44 = B[10];
  assign n_45 = B[10];
  assign n_46 = B[11];
  assign n_47 = B[11];
  assign n_48 = n_0 & n_44;
  assign n_49 = n_48;
  assign n_54 = n_2 & n_24;
  assign n_64 = n_49 & n_54;
  assign n_65 = n_64;
  assign n_126 = n_22 & n_24;
  assign n_127 = n_126;
  assign n_136 = ~n_34;
  assign n_137 = n_136;
  assign n_152 = ~n_65;
  assign n_153 = n_152;
  assign n_156 = n_6 & n_26;
  assign n_157 = n_156;
  assign n_214 = ~n_22;
  assign n_215 = n_214;
  assign n_270 = n_215 & n_4;
  assign n_280 = n_153;
  assign n_281 = n_280;
  assign n_380 = n_22 & n_28;
  MUX2X1 tmp78(.Y(n_392), .A(n_137), .B(n_270), .S(n_127));
  assign n_393 = n_392;
  assign n_532 = n_18;
  assign n_540 = n_20 & n_30;
  assign n_548 = n_22 & n_30;
  assign n_620 = n_157 & n_532;
  assign n_621 = n_620;
  assign n_626 = n_380 & n_540;
  assign n_627 = n_626;
  assign n_648 = n_4 & n_32;
  assign n_649 = n_648;
  assign n_692 = n_16 & n_32;
  assign n_700 = n_18 & n_32;
  assign n_704 = n_649;
  assign n_706 = n_20 & n_32;
  assign n_707 = n_706;
  assign n_714 = n_22 & n_32;
  assign n_760 = ~n_281;
  assign n_761 = n_760;
  assign n_778 = n_620 & n_692;
  assign n_779 = n_778;
  FAX1 tmp99(.YS(n_786), .YC(n_787), .A(n_626), .B(n_700), .C(n_621));
  FAX1 tmp100(.YS(n_794), .YC(n_795), .A(n_548), .B(n_706), .C(n_627));
  assign n_852 = n_14 & n_34;
  assign n_853 = n_852;
  assign n_858 = n_16 & n_34;
  assign n_866 = n_18 & n_34;
  assign n_874 = n_20 & n_34;
  assign n_880 = n_22 & n_34;
  assign n_932 = n_853;
  assign n_933 = n_932;
  assign n_938 = ~n_778;
  assign n_939 = n_938;
  FAX1 tmp111(.YS(n_946), .YC(n_947), .A(n_786), .B(n_858), .C(n_779));
  FAX1 tmp112(.YS(n_952), .YC(n_953), .A(n_794), .B(n_866), .C(n_787));
  FAX1 tmp113(.YS(n_960), .YC(n_961), .A(n_714), .B(n_874), .C(n_795));
  assign n_994 = ~n_761;
  assign n_995 = n_994;
  assign n_1010 = n_12 & n_36;
  assign n_1018 = n_14 & n_36;
  assign n_1026 = n_16 & n_36;
  assign n_1032 = n_18 & n_36;
  assign n_1040 = n_20 & n_36;
  assign n_1048 = n_22 & n_36;
  assign n_1054 = n_995;
  FAX1 tmp123(.YS(n_1098), .YC(n_1099), .A(n_938), .B(n_1010), .C(n_933));
  FAX1 tmp124(.YS(n_1104), .YC(n_1105), .A(n_946), .B(n_1018), .C(n_939));
  FAX1 tmp125(.YS(n_1112), .YC(n_1113), .A(n_952), .B(n_1026), .C(n_947));
  FAX1 tmp126(.YS(n_1120), .YC(n_1121), .A(n_960), .B(n_1032), .C(n_953));
  FAX1 tmp127(.YS(n_1126), .YC(n_1127), .A(n_880), .B(n_1040), .C(n_961));
  assign n_1176 = ~n_281;
  assign n_1178 = n_12 & n_38;
  assign n_1184 = n_14 & n_38;
  assign n_1192 = n_16 & n_38;
  assign n_1200 = n_18 & n_38;
  assign n_1206 = n_20 & n_38;
  assign n_1214 = n_22 & n_38;
  assign n_1258 = n_1098;
  assign n_1259 = n_1258;
  FAX1 tmp137(.YS(n_1264), .YC(n_1265), .A(n_1104), .B(n_1178), .C(n_1099));
  FAX1 tmp138(.YS(n_1272), .YC(n_1273), .A(n_1112), .B(n_1184), .C(n_1105));
  FAX1 tmp139(.YS(n_1278), .YC(n_1279), .A(n_1120), .B(n_1192), .C(n_1113));
  FAX1 tmp140(.YS(n_1286), .YC(n_1287), .A(n_1126), .B(n_1200), .C(n_1121));
  FAX1 tmp141(.YS(n_1294), .YC(n_1295), .A(n_1048), .B(n_1206), .C(n_1127));
  assign n_1336 = n_10 & n_40;
  assign n_1344 = n_12 & n_40;
  assign n_1352 = n_14 & n_40;
  assign n_1358 = n_16 & n_40;
  assign n_1366 = n_18 & n_40;
  assign n_1374 = n_20 & n_40;
  assign n_1380 = n_22 & n_40;
  assign n_1388 = ~n_393;
  FAX1 tmp150(.YS(n_1424), .YC(n_1425), .A(n_1264), .B(n_1336), .C(n_1259));
  FAX1 tmp151(.YS(n_1432), .YC(n_1433), .A(n_1272), .B(n_1344), .C(n_1265));
  FAX1 tmp152(.YS(n_1438), .YC(n_1439), .A(n_1278), .B(n_1352), .C(n_1273));
  FAX1 tmp153(.YS(n_1446), .YC(n_1447), .A(n_1286), .B(n_1358), .C(n_1279));
  FAX1 tmp154(.YS(n_1452), .YC(n_1453), .A(n_1294), .B(n_1366), .C(n_1287));
  FAX1 tmp155(.YS(n_1460), .YC(n_1461), .A(n_1214), .B(n_1374), .C(n_1295));
  assign n_1490 = n_6 & n_648;
  assign n_1491 = n_1490;
  assign n_1504 = n_10 & n_42;
  assign n_1510 = n_12 & n_42;
  assign n_1518 = n_14 & n_42;
  assign n_1526 = n_16 & n_42;
  assign n_1532 = n_18 & n_42;
  assign n_1540 = n_20 & n_42;
  assign n_1548 = n_22 & n_42;
  HAX1 tmp165(.YS(n_1584), .YC(n_1585), .A(n_1424), .B(n_1526));
  FAX1 tmp166(.YS(n_1590), .YC(n_1591), .A(n_1432), .B(n_1504), .C(n_1425));
  FAX1 tmp167(.YS(n_1598), .YC(n_1599), .A(n_1438), .B(n_1510), .C(n_1433));
  FAX1 tmp168(.YS(n_1604), .YC(n_1605), .A(n_1446), .B(n_1518), .C(n_1439));
  FAX1 tmp169(.YS(n_1612), .YC(n_1613), .A(n_1452), .B(n_1526), .C(n_1447));
  FAX1 tmp170(.YS(n_1620), .YC(n_1621), .A(n_1460), .B(n_1532), .C(n_1453));
  FAX1 tmp171(.YS(n_1626), .YC(n_1627), .A(n_1380), .B(n_1540), .C(n_1461));
  assign n_1642 = n_2 & n_44;
  assign n_1656 = n_6 & n_44;
  assign n_1662 = n_8 & n_44;
  assign n_1670 = n_10 & n_44;
  assign n_1678 = n_12 & n_44;
  assign n_1684 = n_14 & n_44;
  assign n_1692 = n_16 & n_44;
  assign n_1700 = n_18 & n_44;
  assign n_1706 = n_20 & n_44;
  assign n_1714 = n_22 & n_44;
  assign n_1742 = n_1584 | n_1656;
  assign n_1743 = n_1742;
  FAX1 tmp184(.YS(n_1750), .YC(n_1751), .A(n_1590), .B(n_1662), .C(n_1585));
  FAX1 tmp185(.YS(n_1758), .YC(n_1759), .A(n_1598), .B(n_1670), .C(n_1591));
  FAX1 tmp186(.YS(n_1764), .YC(n_1765), .A(n_1604), .B(n_1678), .C(n_1599));
  FAX1 tmp187(.YS(n_1772), .YC(n_1773), .A(n_1612), .B(n_1684), .C(n_1605));
  FAX1 tmp188(.YS(n_1778), .YC(n_1779), .A(n_1620), .B(n_1692), .C(n_1613));
  FAX1 tmp189(.YS(n_1786), .YC(n_1787), .A(n_1626), .B(n_1700), .C(n_1621));
  FAX1 tmp190(.YS(n_1794), .YC(n_1795), .A(n_1548), .B(n_1706), .C(n_1627));
  assign n_1822 = n_6 & n_46;
  assign n_1830 = n_8 & n_46;
  assign n_1836 = n_10 & n_46;
  assign n_1837 = n_1836;
  assign n_1844 = n_12 & n_46;
  assign n_1852 = n_14 & n_46;
  assign n_1858 = n_16 & n_46;
  assign n_1866 = n_18 & n_46;
  assign n_1874 = n_20 & n_46;
  assign n_1880 = n_22 & n_46;
  assign n_1902 = n_707;
  assign n_1903 = n_1902;
  FAX1 tmp203(.YS(n_1910), .YC(n_1911), .A(n_779), .B(n_1822), .C(n_1743));
  FAX1 tmp204(.YS(n_1916), .YC(n_1917), .A(n_1758), .B(n_1830), .C(n_1751));
  FAX1 tmp205(.YS(n_1924), .YC(n_1925), .A(n_1764), .B(n_1836), .C(n_1759));
  FAX1 tmp206(.YS(n_1932), .YC(n_1933), .A(n_1772), .B(n_1844), .C(n_1765));
  FAX1 tmp207(.YS(n_1938), .YC(n_1939), .A(n_1778), .B(n_1852), .C(n_1773));
  FAX1 tmp208(.YS(n_1946), .YC(n_1947), .A(n_1786), .B(n_1858), .C(n_1779));
  FAX1 tmp209(.YS(n_1952), .YC(n_1953), .A(n_1794), .B(n_1866), .C(n_1787));
  FAX1 tmp210(.YS(n_1960), .YC(n_1961), .A(n_1714), .B(n_1874), .C(n_1795));
  assign n_1974 = ~n_1902;
  HAX1 tmp212(.YS(n_1982), .YC(n_1983), .A(n_1910), .B(n_1903));
  FAX1 tmp213(.YS(n_1990), .YC(n_1991), .A(n_1916), .B(n_1911), .C(n_1983));
  FAX1 tmp214(.YS(n_1996), .YC(n_1997), .A(n_1924), .B(n_1917), .C(n_1991));
  FAX1 tmp215(.YS(n_2004), .YC(n_2005), .A(n_1932), .B(n_1925), .C(n_1997));
  FAX1 tmp216(.YS(n_2010), .YC(n_2011), .A(n_1938), .B(n_1933), .C(n_2005));
  FAX1 tmp217(.YS(n_2018), .YC(n_2019), .A(n_1946), .B(n_1939), .C(n_2011));
  FAX1 tmp218(.YS(n_2026), .YC(n_2027), .A(n_1952), .B(n_1947), .C(n_2019));
  FAX1 tmp219(.YS(n_2032), .YC(n_2033), .A(n_1960), .B(n_1953), .C(n_2027));
  FAX1 tmp220(.YS(n_2040), .YC(n_2041), .A(n_1880), .B(n_1961), .C(n_2033));
  assign O[0] = n_48;
  assign O[1] = n_12;
  assign O[2] = n_22;
  assign O[3] = n_704;
  assign O[4] = n_1933;
  assign O[5] = n_1642;
  assign O[6] = n_1054;
  assign O[7] = n_532;
  assign O[8] = n_1388;
  assign O[9] = n_1526;
  assign O[10] = n_1491;
  assign O[11] = n_1176;
  assign O[12] = n_1837;
  assign O[13] = n_1974;
  assign O[14] = n_1982;
  assign O[15] = n_1990;
  assign O[16] = n_1996;
  assign O[17] = n_2004;
  assign O[18] = n_2010;
  assign O[19] = n_2018;
  assign O[20] = n_2026;
  assign O[21] = n_2032;
  assign O[22] = n_2040;
  assign O[23] = n_2041;
endmodule


// internal reference: cgp-compare17.12.mul12u_pwr_0_427_mae_00_0729

