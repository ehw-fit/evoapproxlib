/***
* This code is a part of EvoApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under The MIT License.
* When used, please cite the following article(s): V. Mrazek, R. Hrbacek, Z. Vasicek and L. Sekanina, "EvoApprox8b: Library of approximate adders and multipliers for circuit design and benchmarking of approximation methods". Design, Automation & Test in Europe Conference & Exhibition (DATE), 2017, Lausanne, 2017, pp. 258-261. doi: 10.23919/DATE.2017.7926993 
* This file contains a circuit from a sub-set of pareto optimal circuits with respect to the pwr and mre parameters
***/
// MAE% = 0.059 %
// MAE = 38 
// WCE% = 0.45 %
// WCE = 292 
// WCRE% = 43.56 %
// EP% = 69.26 %
// MRE% = 0.80 %
// MSE = 3147 
// PDK45_PWR = 0.304 mW
// PDK45_AREA = 590.4 um2
// PDK45_DELAY = 1.13 ns

module mul8u_ZFB (
    A,
    B,
    O
);

input [7:0] A;
input [7:0] B;
output [15:0] O;

wire sig_16,sig_17,sig_18,sig_19,sig_20,sig_21,sig_22,sig_23,sig_24,sig_25,sig_26,sig_27,sig_28,sig_29,sig_30,sig_31,sig_32,sig_33,sig_34,sig_35;
wire sig_36,sig_37,sig_38,sig_39,sig_40,sig_41,sig_42,sig_43,sig_44,sig_45,sig_46,sig_47,sig_48,sig_49,sig_50,sig_51,sig_52,sig_53,sig_54,sig_55;
wire sig_56,sig_57,sig_58,sig_59,sig_60,sig_61,sig_62,sig_63,sig_64,sig_65,sig_66,sig_67,sig_68,sig_69,sig_70,sig_71,sig_72,sig_73,sig_74,sig_75;
wire sig_76,sig_77,sig_78,sig_79,sig_80,sig_82,sig_85,sig_87,sig_90,sig_92,sig_95,sig_97,sig_100,sig_102,sig_103,sig_104,sig_105,sig_106,sig_107,sig_108;
wire sig_109,sig_110,sig_111,sig_112,sig_113,sig_114,sig_116,sig_117,sig_119,sig_121,sig_122,sig_123,sig_124,sig_125,sig_126,sig_127,sig_128,sig_129,sig_130,sig_131;
wire sig_132,sig_133,sig_134,sig_135,sig_136,sig_137,sig_138,sig_139,sig_140,sig_141,sig_142,sig_143,sig_144,sig_145,sig_146,sig_147,sig_153,sig_158,sig_163,sig_166;
wire sig_168,sig_170,sig_171,sig_172,sig_173,sig_174,sig_175,sig_176,sig_177,sig_178,sig_179,sig_180,sig_181,sig_182,sig_183,sig_184,sig_185,sig_187,sig_188,sig_189;
wire sig_190,sig_191,sig_192,sig_193,sig_194,sig_195,sig_196,sig_197,sig_198,sig_199,sig_200,sig_201,sig_202,sig_203,sig_204,sig_205,sig_206,sig_207,sig_208,sig_209;
wire sig_210,sig_211,sig_212,sig_213,sig_214,sig_215,sig_216,sig_217,sig_218,sig_230,sig_231,sig_233,sig_234,sig_235,sig_236,sig_237,sig_238,sig_239,sig_240,sig_241;
wire sig_242,sig_243,sig_244,sig_245,sig_246,sig_247,sig_248,sig_249,sig_250,sig_251,sig_252,sig_253,sig_254,sig_255,sig_256,sig_262,sig_264,sig_268,sig_269,sig_270;
wire sig_271,sig_272,sig_273,sig_274,sig_275,sig_276,sig_277,sig_278,sig_279,sig_280,sig_281,sig_282,sig_283,sig_284,sig_285,sig_286,sig_287,sig_288,sig_289,sig_290;
wire sig_291,sig_292,sig_293,sig_294,sig_295,sig_296,sig_297,sig_298,sig_299,sig_305,sig_306,sig_307,sig_308,sig_309,sig_310,sig_311,sig_312,sig_313,sig_314,sig_315;
wire sig_316,sig_317,sig_318,sig_319,sig_353,sig_356,sig_358,sig_363,sig_367,sig_368,sig_370,sig_372,sig_374,sig_378,sig_382,sig_383,sig_389,sig_390,sig_391,sig_401;
wire sig_402,sig_404,sig_405,sig_407,sig_409,sig_411,sig_425,sig_432,sig_434,sig_435,sig_437,sig_448,sig_451,sig_452,sig_456,sig_457,sig_463,sig_464,sig_498,sig_499;
wire sig_500,sig_501,sig_502,sig_503,sig_504,sig_505;

assign sig_16 = B[0] & A[0];
assign sig_17 = B[1] & A[0];
assign sig_18 = B[2] & A[0];
assign sig_19 = B[3] & A[0];
assign sig_20 = B[4] & A[0];
assign sig_21 = B[5] & A[0];
assign sig_22 = B[6] & A[0];
assign sig_23 = B[7] & A[0];
assign sig_24 = B[0] & A[1];
assign sig_25 = B[1] & A[1];
assign sig_26 = B[2] & A[1];
assign sig_27 = B[3] & A[1];
assign sig_28 = B[4] & A[1];
assign sig_29 = B[5] & A[1];
assign sig_30 = B[6] & A[1];
assign sig_31 = B[7] & A[1];
assign sig_32 = B[0] & A[2];
assign sig_33 = B[1] & A[2];
assign sig_34 = B[2] & A[2];
assign sig_35 = B[3] & A[2];
assign sig_36 = B[4] & A[2];
assign sig_37 = B[5] & A[2];
assign sig_38 = B[6] & A[2];
assign sig_39 = B[7] & A[2];
assign sig_40 = B[0] & A[3];
assign sig_41 = B[1] & A[3];
assign sig_42 = B[2] & A[3];
assign sig_43 = B[3] & A[3];
assign sig_44 = B[4] & A[3];
assign sig_45 = B[5] & A[3];
assign sig_46 = B[6] & A[3];
assign sig_47 = B[7] & A[3];
assign sig_48 = B[0] & A[4];
assign sig_49 = B[1] & A[4];
assign sig_50 = B[2] & A[4];
assign sig_51 = B[3] & A[4];
assign sig_52 = B[4] & A[4];
assign sig_53 = B[5] & A[4];
assign sig_54 = B[6] & A[4];
assign sig_55 = B[7] & A[4];
assign sig_56 = B[0] & A[5];
assign sig_57 = B[1] & A[5];
assign sig_58 = B[2] & A[5];
assign sig_59 = B[3] & A[5];
assign sig_60 = B[4] & A[5];
assign sig_61 = B[5] & A[5];
assign sig_62 = B[6] & A[5];
assign sig_63 = B[7] & A[5];
assign sig_64 = B[0] & A[6];
assign sig_65 = B[1] & A[6];
assign sig_66 = B[2] & A[6];
assign sig_67 = B[3] & A[6];
assign sig_68 = B[4] & A[6];
assign sig_69 = B[5] & A[6];
assign sig_70 = B[6] & A[6];
assign sig_71 = B[7] & A[6];
assign sig_72 = B[0] & A[7];
assign sig_73 = B[1] & A[7];
assign sig_74 = B[2] & A[7];
assign sig_75 = B[3] & A[7];
assign sig_76 = B[4] & A[7];
assign sig_77 = B[5] & A[7];
assign sig_78 = B[6] & A[7];
assign sig_79 = B[7] & A[7];
assign sig_80 = sig_17 | sig_24;
assign sig_82 = sig_18 | sig_25;
assign sig_85 = sig_82 | sig_32;
assign sig_87 = sig_19 | sig_26;
assign sig_90 = sig_87 | sig_33;
assign sig_92 = sig_20 | sig_27;
assign sig_95 = sig_92 | sig_34;
assign sig_97 = sig_21 | sig_28;
assign sig_100 = sig_97 | sig_35;
assign sig_102 = sig_22 | sig_29;
assign sig_103 = sig_22 & sig_29;
assign sig_104 = sig_102 & sig_36;
assign sig_105 = sig_102 | sig_36;
assign sig_106 = sig_103 | sig_104;
assign sig_107 = sig_23 ^ sig_30;
assign sig_108 = sig_23 & sig_30;
assign sig_109 = sig_107 & sig_37;
assign sig_110 = sig_107 ^ sig_37;
assign sig_111 = sig_108 | sig_109;
assign sig_112 = sig_31 & sig_38;
assign sig_113 = sig_31 ^ sig_38;
assign sig_114 = sig_41 | sig_48;
assign sig_116 = sig_42 | sig_49;
assign sig_117 = sig_42 & B[5];
assign sig_119 = sig_116 | sig_56;
assign sig_121 = sig_43 ^ sig_50;
assign sig_122 = sig_43 & sig_50;
assign sig_123 = sig_121 & sig_57;
assign sig_124 = sig_121 ^ sig_57;
assign sig_125 = sig_122 | sig_123;
assign sig_126 = sig_44 ^ sig_51;
assign sig_127 = sig_44 & sig_51;
assign sig_128 = sig_126 & sig_58;
assign sig_129 = sig_126 ^ sig_58;
assign sig_130 = sig_127 | sig_128;
assign sig_131 = sig_45 ^ sig_52;
assign sig_132 = sig_45 & sig_52;
assign sig_133 = sig_131 & sig_59;
assign sig_134 = sig_131 ^ sig_59;
assign sig_135 = sig_132 | sig_133;
assign sig_136 = sig_46 ^ sig_53;
assign sig_137 = sig_46 & sig_53;
assign sig_138 = sig_136 & sig_60;
assign sig_139 = sig_136 ^ sig_60;
assign sig_140 = sig_137 | sig_138;
assign sig_141 = sig_47 ^ sig_54;
assign sig_142 = sig_47 & sig_54;
assign sig_143 = sig_141 & sig_61;
assign sig_144 = sig_141 ^ sig_61;
assign sig_145 = sig_142 | sig_143;
assign sig_146 = sig_55 & sig_62;
assign sig_147 = sig_55 ^ sig_62;
assign sig_153 = sig_90 | sig_40;
assign sig_158 = sig_95 | sig_114;
assign sig_163 = sig_100 | sig_119;
assign sig_166 = sig_105 & sig_124;
assign sig_168 = sig_105 | sig_124;
assign sig_170 = sig_110 ^ sig_106;
assign sig_171 = sig_110 & sig_106;
assign sig_172 = sig_170 & sig_129;
assign sig_173 = sig_170 ^ sig_129;
assign sig_174 = sig_171 | sig_172;
assign sig_175 = sig_113 ^ sig_111;
assign sig_176 = sig_113 & sig_111;
assign sig_177 = sig_175 & sig_134;
assign sig_178 = sig_175 ^ sig_134;
assign sig_179 = sig_176 | sig_177;
assign sig_180 = sig_39 ^ sig_112;
assign sig_181 = B[6] & sig_112;
assign sig_182 = sig_180 & sig_139;
assign sig_183 = sig_180 ^ sig_139;
assign sig_184 = sig_181 | sig_182;
assign sig_185 = sig_117 | sig_64;
assign sig_187 = sig_125 ^ sig_65;
assign sig_188 = sig_125 & sig_65;
assign sig_189 = sig_187 & sig_72;
assign sig_190 = sig_187 | sig_72;
assign sig_191 = sig_188 | sig_189;
assign sig_192 = sig_130 ^ sig_66;
assign sig_193 = sig_130 & sig_66;
assign sig_194 = sig_192 & sig_73;
assign sig_195 = sig_192 ^ sig_73;
assign sig_196 = sig_193 | sig_194;
assign sig_197 = sig_135 ^ sig_67;
assign sig_198 = sig_135 & sig_67;
assign sig_199 = sig_197 & sig_74;
assign sig_200 = sig_197 ^ sig_74;
assign sig_201 = sig_198 | sig_199;
assign sig_202 = sig_140 ^ sig_68;
assign sig_203 = sig_140 & sig_68;
assign sig_204 = sig_202 & sig_75;
assign sig_205 = sig_202 ^ sig_75;
assign sig_206 = sig_203 | sig_204;
assign sig_207 = sig_145 ^ sig_69;
assign sig_208 = sig_145 & sig_69;
assign sig_209 = sig_207 & sig_76;
assign sig_210 = sig_207 ^ sig_76;
assign sig_211 = sig_208 | sig_209;
assign sig_212 = sig_146 ^ sig_70;
assign sig_213 = sig_146 & sig_70;
assign sig_214 = sig_212 & sig_77;
assign sig_215 = sig_212 ^ sig_77;
assign sig_216 = sig_213 | sig_214;
assign sig_217 = sig_71 & A[7];
assign sig_218 = sig_71 ^ sig_78;
assign sig_230 = sig_188 & sig_185;
assign sig_231 = sig_168 | sig_185;
assign sig_233 = sig_173 ^ sig_166;
assign sig_234 = sig_173 & sig_166;
assign sig_235 = sig_233 & sig_190;
assign sig_236 = sig_233 ^ sig_190;
assign sig_237 = sig_234 | sig_235;
assign sig_238 = sig_178 ^ sig_174;
assign sig_239 = sig_178 & sig_174;
assign sig_240 = sig_238 & sig_195;
assign sig_241 = sig_238 ^ sig_195;
assign sig_242 = sig_239 | sig_240;
assign sig_243 = sig_183 ^ sig_179;
assign sig_244 = sig_183 & sig_179;
assign sig_245 = sig_243 & sig_200;
assign sig_246 = sig_243 ^ sig_200;
assign sig_247 = sig_244 | sig_245;
assign sig_248 = sig_144 ^ sig_184;
assign sig_249 = sig_144 & sig_184;
assign sig_250 = sig_248 & sig_205;
assign sig_251 = sig_248 ^ sig_205;
assign sig_252 = sig_249 | sig_250;
assign sig_253 = sig_147 & sig_210;
assign sig_254 = sig_147 ^ sig_210;
assign sig_255 = sig_63 & sig_215;
assign sig_256 = sig_63 ^ sig_215;
assign sig_262 = A[2] & sig_235;
assign sig_264 = A[1] & sig_230;
assign sig_268 = sig_241 ^ sig_237;
assign sig_269 = sig_241 & sig_237;
assign sig_270 = sig_268 & sig_191;
assign sig_271 = sig_268 ^ sig_191;
assign sig_272 = sig_269 | sig_270;
assign sig_273 = sig_246 ^ sig_242;
assign sig_274 = sig_246 & sig_242;
assign sig_275 = sig_273 & sig_196;
assign sig_276 = sig_273 ^ sig_196;
assign sig_277 = sig_274 | sig_275;
assign sig_278 = sig_251 ^ sig_247;
assign sig_279 = sig_251 & sig_247;
assign sig_280 = sig_278 & sig_201;
assign sig_281 = sig_278 ^ sig_201;
assign sig_282 = sig_279 | sig_280;
assign sig_283 = sig_254 ^ sig_252;
assign sig_284 = sig_254 & sig_252;
assign sig_285 = sig_283 & sig_206;
assign sig_286 = sig_283 ^ sig_206;
assign sig_287 = sig_284 | sig_285;
assign sig_288 = sig_256 ^ sig_253;
assign sig_289 = sig_256 & sig_253;
assign sig_290 = sig_288 & sig_211;
assign sig_291 = sig_288 ^ sig_211;
assign sig_292 = sig_289 | sig_290;
assign sig_293 = sig_218 ^ sig_255;
assign sig_294 = sig_218 & sig_255;
assign sig_295 = sig_293 & sig_216;
assign sig_296 = sig_293 ^ sig_216;
assign sig_297 = sig_294 | sig_295;
assign sig_298 = B[6] & sig_217;
assign sig_299 = sig_79 ^ sig_298;
assign sig_305 = sig_236 & sig_262;
assign sig_306 = sig_271 ^ sig_264;
assign sig_307 = sig_271 & sig_264;
assign sig_308 = sig_276 ^ sig_272;
assign sig_309 = sig_276 & sig_272;
assign sig_310 = sig_281 ^ sig_277;
assign sig_311 = sig_281 & sig_277;
assign sig_312 = sig_286 ^ sig_282;
assign sig_313 = sig_286 & sig_282;
assign sig_314 = sig_291 ^ sig_287;
assign sig_315 = sig_291 & sig_287;
assign sig_316 = sig_296 ^ sig_292;
assign sig_317 = sig_296 & sig_292;
assign sig_318 = sig_299 ^ sig_297;
assign sig_319 = sig_299 & sig_297;
assign sig_353 = sig_308 & sig_307;
assign sig_356 = sig_353 | sig_309;
assign sig_358 = sig_310 & sig_308;
assign sig_363 = sig_358 & sig_356;
assign sig_367 = sig_310 & sig_309;
assign sig_368 = sig_311 | sig_367;
assign sig_370 = sig_305 | sig_363;
assign sig_372 = sig_368 | sig_370;
assign sig_374 = sig_307 & B[1];
assign sig_378 = sig_312 & sig_363;
assign sig_382 = sig_374 & sig_358;
assign sig_383 = sig_312 & sig_368;
assign sig_389 = sig_383 | sig_378;
assign sig_390 = sig_313 | sig_389;
assign sig_391 = sig_314 & sig_312;
assign sig_401 = sig_391 & sig_382;
assign sig_402 = sig_391 & sig_368;
assign sig_404 = sig_314 & sig_313;
assign sig_405 = sig_315 | sig_404;
assign sig_407 = sig_401 | sig_404;
assign sig_409 = sig_405 | sig_402;
assign sig_411 = sig_409 | sig_407;
assign sig_425 = sig_316 & sig_409;
assign sig_432 = sig_316 & sig_407;
assign sig_434 = sig_425 | sig_432;
assign sig_435 = sig_317 | sig_434;
assign sig_437 = sig_318 & sig_316;
assign sig_448 = sig_437 & sig_391;
assign sig_451 = sig_448 & sig_382;
assign sig_452 = sig_437 & sig_409;
assign sig_456 = sig_318 & sig_317;
assign sig_457 = sig_319 | sig_456;
assign sig_463 = sig_452 | sig_457;
assign sig_464 = sig_451 | sig_463;
assign sig_498 = sig_306 ^ sig_305;
assign sig_499 = sig_308 ^ sig_307;
assign sig_500 = sig_310 ^ sig_356;
assign sig_501 = sig_312 ^ sig_372;
assign sig_502 = sig_314 ^ sig_390;
assign sig_503 = sig_316 ^ sig_411;
assign sig_504 = sig_318 ^ sig_435;
assign sig_505 = sig_298 | sig_464;

assign O[15] = sig_505;
assign O[14] = sig_504;
assign O[13] = sig_503;
assign O[12] = sig_502;
assign O[11] = sig_501;
assign O[10] = sig_500;
assign O[9] = sig_499;
assign O[8] = sig_498;
assign O[7] = sig_236;
assign O[6] = sig_231;
assign O[5] = sig_163;
assign O[4] = sig_158;
assign O[3] = sig_153;
assign O[2] = sig_85;
assign O[1] = sig_80;
assign O[0] = sig_16;

endmodule


