/***
* This code is a part of ApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under a XXXX public license.
* When used, please cite the following article: tbd 
* This file is pareto optimal sub-set in the pdk45_pwr and mae% parameters
***/

module mul12u_pwr_0_709_mae_00_0109(A, B, O);
  input [11:0] A, B;
  output [23:0] O;
  wire n_1198, n_1199, n_1190, n_1191, n_1619, n_1618, n_1754, n_1755, n_1204, n_1612;
  wire n_1682, n_706, n_488, n_489, n_1103, n_1102, n_1109, n_1108, n_1295, n_1294;
  wire n_1862, n_1863, n_1868, n_1869, n_724, n_2034, n_2035, n_1613, n_552, n_654;
  wire n_558, n_1408, n_1409, n_1033, n_1032, n_832, n_1976, n_424, n_1038, n_1402;
  wire n_1403, n_348, n_18, n_19, n_16, n_17, n_14, n_15, n_12, n_13;
  wire n_10, n_11, n_1729, n_334, n_336, n_337, n_1536, n_1537, n_1530, n_1242;
  wire n_1243, n_1248, n_1249, n_906, n_1082, n_904, n_86, n_1912, n_1664, n_1985;
  wire n_1984, n_564, n_162, n_1581, n_264, n_1580, n_794, n_762, n_415, n_414;
  wire n_1365, n_942, n_412, n_418, n_948, n_45, n_44, n_47, n_46, n_41;
  wire n_40, n_43, n_42, n_864, n_1958, n_1959, n_49, n_48, n_1895, n_1894;
  wire n_1562, n_468, n_1446, n_1440, n_1441, n_1569, n_1568, n_1626, n_1627, n_1185;
  wire n_1184, n_1747, n_1746, n_1217, n_1216, n_1211, n_1210, n_1741, n_1740, n_8;
  wire n_9, n_1875, n_1874, n_182, n_634, n_188, n_224, n_225, n_2023, n_2022;
  wire n_1452, n_2029, n_2028, n_648, n_642, n_820, n_352, n_826, n_1554, n_1555;
  wire n_1000, n_1001, n_730, n_738, n_739, n_1638, n_1255, n_1254, n_1095, n_1094;
  wire n_916, n_910, n_858, n_78, n_1906, n_1901, n_1900, n_72, n_73, n_1415;
  wire n_1414, n_1798, n_1799, n_1792, n_1172, n_1173, n_1178, n_1179, n_1772, n_1773;
  wire n_1676, n_1778, n_1670, n_1831, n_1830, n_1837, n_1836, n_578, n_570, n_176;
  wire n_177, n_253, n_252, n_707, n_258, n_316, n_852, n_1364, n_2016, n_2017;
  wire n_675, n_674, n_770, n_776, n_404, n_954, n_1428, n_1429, n_1356, n_1357;
  wire n_1350, n_1351, n_1420, n_1421, n_30, n_31, n_32, n_33, n_34, n_35;
  wire n_36, n_37, n_38, n_39, n_1952, n_1453, n_494, n_1633, n_1632, n_1639;
  wire n_782, n_922, n_1222, n_1223, n_928, n_1734, n_1735, n_1044, n_788, n_1644;
  wire n_1645, n_1127, n_1126, n_1120, n_1842, n_1843, n_1848, n_1849, n_198, n_628;
  wire n_194, n_622, n_532, n_109, n_108, n_1965, n_1964, n_104, n_1019, n_1018;
  wire n_1549, n_1548, n_1543, n_1542, n_692, n_698, n_2041, n_2040, n_744, n_1045;
  wire n_1268, n_1269, n_1262, n_1263, n_846, n_840, n_960, n_67, n_66, n_1460;
  wire n_1466, n_1671, n_1787, n_1786, n_1167, n_1166, n_4, n_5, n_6, n_7;
  wire n_0, n_1, n_2, n_3, n_1767, n_1766, n_1761, n_1760, n_1600, n_1601;
  wire n_1606, n_1607, n_540, n_546, n_1114, n_1115, n_1286, n_1280, n_1281, n_145;
  wire n_144, n_202, n_2009, n_718, n_2008, n_712, n_392, n_393, n_398, n_2002;
  wire n_2003, n_1024, n_1025, n_1435, n_1434, n_1083, n_23, n_22, n_21, n_20;
  wire n_27, n_26, n_25, n_24, n_29, n_28, n_1970, n_1971, n_890, n_897;
  wire n_896, n_482, n_328, n_1237, n_1236, n_1231, n_1230, n_936, n_1728, n_1926;
  wire n_1158, n_1159, n_1651, n_1650, n_1152, n_1153, n_1659, n_1658, n_1996, n_1997;
  wire n_1990, n_1991, n_1857, n_1856, n_610, n_616, n_340, n_118, n_808, n_500;
  wire n_270, n_273, n_272, n_1574, n_686, n_680, n_800, n_884, n_1977, n_750;
  wire n_203, n_756, n_1370, n_1371, n_1275, n_1274, n_872, n_1888, n_1889, n_1920;
  wire n_878, n_1880, n_1881, n_58, n_59, n_52, n_53, n_54, n_476, n_1472;
  wire n_1479, n_1478;
  assign n_0 = A[0];
  assign n_1 = A[0];
  assign n_2 = A[1];
  assign n_3 = A[1];
  assign n_4 = A[2];
  assign n_5 = A[2];
  assign n_6 = A[3];
  assign n_7 = A[3];
  assign n_8 = A[4];
  assign n_9 = A[4];
  assign n_10 = A[5];
  assign n_11 = A[5];
  assign n_12 = A[6];
  assign n_13 = A[6];
  assign n_14 = A[7];
  assign n_15 = A[7];
  assign n_16 = A[8];
  assign n_17 = A[8];
  assign n_18 = A[9];
  assign n_19 = A[9];
  assign n_20 = A[10];
  assign n_21 = A[10];
  assign n_22 = A[11];
  assign n_23 = A[11];
  assign n_24 = B[0];
  assign n_25 = B[0];
  assign n_26 = B[1];
  assign n_27 = B[1];
  assign n_28 = B[2];
  assign n_29 = B[2];
  assign n_30 = B[3];
  assign n_31 = B[3];
  assign n_32 = B[4];
  assign n_33 = B[4];
  assign n_34 = B[5];
  assign n_35 = B[5];
  assign n_36 = B[6];
  assign n_37 = B[6];
  assign n_38 = B[7];
  assign n_39 = B[7];
  assign n_40 = B[8];
  assign n_41 = B[8];
  assign n_42 = B[9];
  assign n_43 = B[9];
  assign n_44 = B[10];
  assign n_45 = B[10];
  assign n_46 = B[11];
  assign n_47 = B[11];
  assign n_48 = n_28 & n_12;
  assign n_49 = n_48;
  assign n_52 = ~(n_42 & n_4 & n_46);
  assign n_53 = n_52;
  assign n_54 = ~(n_2 | n_52 | n_42);
  assign n_58 = ~(n_53 | n_42);
  assign n_59 = n_58;
  assign n_66 = ~n_59;
  assign n_67 = n_66;
  assign n_72 = n_2 & n_54;
  assign n_73 = n_72;
  assign n_78 = n_49 & n_32;
  assign n_86 = n_14 & n_16;
  assign n_104 = n_34 & n_78;
  assign n_108 = ~n_73;
  assign n_109 = n_108;
  assign n_118 = n_22 & n_24;
  assign n_144 = n_109;
  assign n_145 = n_144;
  assign n_162 = n_12 & n_26;
  assign n_176 = n_73 & n_54;
  assign n_177 = n_176;
  assign n_182 = n_18 & n_162;
  assign n_188 = n_20 & n_26;
  assign n_194 = n_22 & n_26;
  assign n_198 = ~n_177;
  assign n_202 = ~(n_26 | n_198);
  assign n_203 = n_202;
  assign n_224 = ~n_177;
  assign n_225 = n_224;
  OAI21X1 tmp89(.Y(n_252), .A(n_26), .B(n_66), .C(n_59));
  assign n_253 = n_252;
  assign n_258 = n_18 & n_28;
  assign n_264 = n_20 & n_28;
  assign n_270 = n_22 & n_28;
  assign n_272 = ~n_225;
  assign n_273 = n_272;
  assign n_316 = n_273;
  assign n_328 = n_16 & n_30;
  assign n_334 = n_18 & n_30;
  assign n_336 = ~n_145;
  assign n_337 = n_336;
  assign n_340 = n_20 & n_30;
  assign n_348 = n_22 & n_30;
  assign n_352 = ~n_273;
  OAI21X1 tmp104(.Y(n_392), .A(n_34), .B(n_12), .C(n_203));
  assign n_393 = n_392;
  assign n_398 = n_14 & n_32;
  assign n_404 = n_16 & n_32;
  assign n_412 = n_18 & n_32;
  assign n_414 = ~n_393;
  assign n_415 = n_414;
  assign n_418 = n_20 & n_32;
  assign n_424 = n_22 & n_32;
  assign n_468 = n_12 & n_34;
  assign n_476 = n_14 & n_34;
  assign n_482 = n_16 & n_34;
  assign n_488 = n_18 & n_34;
  assign n_489 = n_488;
  assign n_494 = n_20 & n_34;
  assign n_500 = n_22 & n_34;
  assign n_532 = n_8 & n_36;
  assign n_540 = n_10 & n_36;
  assign n_546 = n_12 & n_36;
  assign n_552 = n_14 & n_36;
  assign n_558 = n_16 & n_36;
  assign n_564 = n_18 & n_36;
  assign n_570 = n_20 & n_36;
  assign n_578 = n_22 & n_36;
  assign n_610 = n_8 & n_38;
  assign n_616 = n_10 & n_38;
  assign n_622 = n_12 & n_38;
  assign n_628 = n_14 & n_38;
  assign n_634 = n_16 & n_38;
  assign n_642 = n_18 & n_38;
  assign n_648 = n_20 & n_38;
  assign n_654 = n_22 & n_38;
  assign n_674 = n_4 & n_40;
  assign n_675 = n_674;
  assign n_680 = n_6 & n_40;
  assign n_686 = n_8 & n_40;
  assign n_692 = n_10 & n_40;
  assign n_698 = n_12 & n_40;
  assign n_706 = n_14 & n_40;
  assign n_707 = n_706;
  assign n_712 = n_16 & n_40;
  assign n_718 = n_18 & n_40;
  assign n_724 = n_20 & n_40;
  assign n_730 = n_22 & n_40;
  assign n_738 = n_0;
  assign n_739 = n_738;
  assign n_744 = ~(n_337 & n_28);
  assign n_750 = n_4 & n_42;
  assign n_756 = n_6 & n_42;
  assign n_762 = n_8 & n_42;
  assign n_770 = n_10 & n_42;
  assign n_776 = n_12 & n_42;
  assign n_782 = n_14 & n_42;
  assign n_788 = n_16 & n_42;
  assign n_794 = n_18 & n_42;
  assign n_800 = n_20 & n_42;
  assign n_808 = n_22 & n_42;
  assign n_820 = n_2 & n_44;
  assign n_826 = n_4 & n_44;
  assign n_832 = n_6 & n_44;
  assign n_840 = n_8 & n_44;
  assign n_846 = n_10 & n_44;
  assign n_852 = n_12 & n_44;
  assign n_858 = n_14 & n_44;
  assign n_864 = n_16 & n_44;
  assign n_872 = n_18 & n_44;
  assign n_878 = n_20 & n_44;
  assign n_884 = n_22 & n_44;
  assign n_890 = n_0 & n_46;
  assign n_896 = n_2 & n_46;
  assign n_897 = n_896;
  assign n_904 = n_4 & n_46;
  assign n_906 = n_253;
  assign n_910 = n_6 & n_46;
  assign n_916 = n_8 & n_46;
  assign n_922 = n_10 & n_46;
  assign n_928 = n_12 & n_46;
  assign n_936 = n_14 & n_46;
  assign n_942 = n_16 & n_46;
  assign n_948 = n_18 & n_46;
  assign n_954 = n_20 & n_46;
  assign n_960 = n_22 & n_46;
  assign n_1000 = n_86 & n_494;
  assign n_1001 = n_1000;
  assign n_1018 = n_104;
  assign n_1019 = n_1018;
  FAX1 tmp190(.YS(n_1024), .YC(n_1025), .A(n_73), .B(n_182), .C(n_67));
  FAX1 tmp191(.YS(n_1032), .YC(n_1033), .A(n_118), .B(n_188), .C(n_258));
  assign n_1038 = n_194 & n_264;
  HAX1 tmp193(.YS(n_1044), .YC(n_1045), .A(n_194), .B(n_264));
  assign n_1082 = n_316;
  assign n_1083 = n_1082;
  FAX1 tmp196(.YS(n_1094), .YC(n_1095), .A(n_328), .B(n_398), .C(n_468));
  FAX1 tmp197(.YS(n_1102), .YC(n_1103), .A(n_334), .B(n_404), .C(n_476));
  FAX1 tmp198(.YS(n_1108), .YC(n_1109), .A(n_340), .B(n_412), .C(n_482));
  FAX1 tmp199(.YS(n_1114), .YC(n_1115), .A(n_348), .B(n_418), .C(n_489));
  assign n_1120 = n_424 & n_494;
  HAX1 tmp201(.YS(n_1126), .YC(n_1127), .A(n_424), .B(n_494));
  FAX1 tmp202(.YS(n_1152), .YC(n_1153), .A(n_532), .B(n_198), .C(n_674));
  FAX1 tmp203(.YS(n_1158), .YC(n_1159), .A(n_540), .B(n_610), .C(n_680));
  FAX1 tmp204(.YS(n_1166), .YC(n_1167), .A(n_546), .B(n_616), .C(n_686));
  FAX1 tmp205(.YS(n_1172), .YC(n_1173), .A(n_552), .B(n_622), .C(n_692));
  FAX1 tmp206(.YS(n_1178), .YC(n_1179), .A(n_558), .B(n_628), .C(n_698));
  FAX1 tmp207(.YS(n_1184), .YC(n_1185), .A(n_564), .B(n_634), .C(n_707));
  FAX1 tmp208(.YS(n_1190), .YC(n_1191), .A(n_570), .B(n_642), .C(n_712));
  FAX1 tmp209(.YS(n_1198), .YC(n_1199), .A(n_578), .B(n_648), .C(n_718));
  assign n_1204 = n_654 & n_724;
  HAX1 tmp211(.YS(n_1210), .YC(n_1211), .A(n_654), .B(n_724));
  assign n_1216 = ~n_744;
  assign n_1217 = n_1216;
  FAX1 tmp214(.YS(n_1222), .YC(n_1223), .A(n_750), .B(n_820), .C(n_890));
  FAX1 tmp215(.YS(n_1230), .YC(n_1231), .A(n_756), .B(n_826), .C(n_897));
  FAX1 tmp216(.YS(n_1236), .YC(n_1237), .A(n_762), .B(n_832), .C(n_904));
  FAX1 tmp217(.YS(n_1242), .YC(n_1243), .A(n_770), .B(n_840), .C(n_910));
  FAX1 tmp218(.YS(n_1248), .YC(n_1249), .A(n_776), .B(n_846), .C(n_916));
  FAX1 tmp219(.YS(n_1254), .YC(n_1255), .A(n_782), .B(n_852), .C(n_922));
  FAX1 tmp220(.YS(n_1262), .YC(n_1263), .A(n_788), .B(n_858), .C(n_928));
  FAX1 tmp221(.YS(n_1268), .YC(n_1269), .A(n_794), .B(n_864), .C(n_936));
  FAX1 tmp222(.YS(n_1274), .YC(n_1275), .A(n_800), .B(n_872), .C(n_942));
  FAX1 tmp223(.YS(n_1280), .YC(n_1281), .A(n_808), .B(n_878), .C(n_948));
  assign n_1286 = n_884 & n_954;
  HAX1 tmp225(.YS(n_1294), .YC(n_1295), .A(n_884), .B(n_954));
  assign n_1350 = n_1024 & n_1019;
  assign n_1351 = n_1350;
  FAX1 tmp228(.YS(n_1356), .YC(n_1357), .A(n_1032), .B(n_1025), .C(n_1094));
  FAX1 tmp229(.YS(n_1364), .YC(n_1365), .A(n_1044), .B(n_1033), .C(n_1102));
  FAX1 tmp230(.YS(n_1370), .YC(n_1371), .A(n_270), .B(n_1038), .C(n_1108));
  MUX2X1 tmp231(.Y(n_1402), .A(n_1083), .B(n_1152), .S(n_675));
  assign n_1403 = n_1402;
  FAX1 tmp233(.YS(n_1408), .YC(n_1409), .A(n_145), .B(n_1158), .C(n_1153));
  FAX1 tmp234(.YS(n_1414), .YC(n_1415), .A(n_1095), .B(n_1166), .C(n_1159));
  FAX1 tmp235(.YS(n_1420), .YC(n_1421), .A(n_1103), .B(n_1172), .C(n_1167));
  FAX1 tmp236(.YS(n_1428), .YC(n_1429), .A(n_1109), .B(n_1178), .C(n_1173));
  FAX1 tmp237(.YS(n_1434), .YC(n_1435), .A(n_1115), .B(n_1184), .C(n_1179));
  FAX1 tmp238(.YS(n_1440), .YC(n_1441), .A(n_1120), .B(n_1190), .C(n_1185));
  assign n_1446 = n_1198 & n_1191;
  HAX1 tmp240(.YS(n_1452), .YC(n_1453), .A(n_1198), .B(n_1191));
  assign n_1460 = n_1210 & n_1199;
  assign n_1466 = n_1210 ^ n_1199;
  assign n_1472 = n_730 & n_1204;
  HAX1 tmp244(.YS(n_1478), .YC(n_1479), .A(n_730), .B(n_1204));
  assign n_1530 = n_2 & n_414;
  FAX1 tmp246(.YS(n_1536), .YC(n_1537), .A(n_1356), .B(n_1351), .C(n_1408));
  FAX1 tmp247(.YS(n_1542), .YC(n_1543), .A(n_1364), .B(n_1357), .C(n_1414));
  FAX1 tmp248(.YS(n_1548), .YC(n_1549), .A(n_1370), .B(n_1365), .C(n_1420));
  FAX1 tmp249(.YS(n_1554), .YC(n_1555), .A(n_1114), .B(n_1371), .C(n_1428));
  assign n_1562 = n_1126 & n_1434;
  HAX1 tmp251(.YS(n_1568), .YC(n_1569), .A(n_1126), .B(n_1434));
  assign n_1574 = n_500 & n_1440;
  HAX1 tmp253(.YS(n_1580), .YC(n_1581), .A(n_500), .B(n_1440));
  HAX1 tmp254(.YS(n_1600), .YC(n_1601), .A(n_1403), .B(n_1222));
  FAX1 tmp255(.YS(n_1606), .YC(n_1607), .A(n_1409), .B(n_1230), .C(n_1223));
  FAX1 tmp256(.YS(n_1612), .YC(n_1613), .A(n_1415), .B(n_1236), .C(n_1231));
  FAX1 tmp257(.YS(n_1618), .YC(n_1619), .A(n_1421), .B(n_1242), .C(n_1237));
  FAX1 tmp258(.YS(n_1626), .YC(n_1627), .A(n_1429), .B(n_1248), .C(n_1243));
  FAX1 tmp259(.YS(n_1632), .YC(n_1633), .A(n_1435), .B(n_1254), .C(n_1249));
  FAX1 tmp260(.YS(n_1638), .YC(n_1639), .A(n_1441), .B(n_1262), .C(n_1255));
  FAX1 tmp261(.YS(n_1644), .YC(n_1645), .A(n_1446), .B(n_1268), .C(n_1263));
  FAX1 tmp262(.YS(n_1650), .YC(n_1651), .A(n_1460), .B(n_1274), .C(n_1269));
  FAX1 tmp263(.YS(n_1658), .YC(n_1659), .A(n_1472), .B(n_1280), .C(n_1275));
  assign n_1664 = n_1294 & n_1281;
  HAX1 tmp265(.YS(n_1670), .YC(n_1671), .A(n_1294), .B(n_1281));
  assign n_1676 = n_960 & n_1286;
  assign n_1682 = n_960 ^ n_1286;
  assign n_1728 = n_1530;
  assign n_1729 = n_1728;
  FAX1 tmp270(.YS(n_1734), .YC(n_1735), .A(n_1536), .B(n_1728), .C(n_1600));
  FAX1 tmp271(.YS(n_1740), .YC(n_1741), .A(n_1542), .B(n_1537), .C(n_1606));
  FAX1 tmp272(.YS(n_1746), .YC(n_1747), .A(n_1548), .B(n_1543), .C(n_1612));
  FAX1 tmp273(.YS(n_1754), .YC(n_1755), .A(n_1554), .B(n_1549), .C(n_1618));
  FAX1 tmp274(.YS(n_1760), .YC(n_1761), .A(n_1568), .B(n_1555), .C(n_1626));
  FAX1 tmp275(.YS(n_1766), .YC(n_1767), .A(n_1580), .B(n_1562), .C(n_1632));
  FAX1 tmp276(.YS(n_1772), .YC(n_1773), .A(n_1452), .B(n_1574), .C(n_1638));
  assign n_1778 = n_1466 & n_1644;
  HAX1 tmp278(.YS(n_1786), .YC(n_1787), .A(n_1466), .B(n_1644));
  assign n_1792 = n_1478 & n_1650;
  HAX1 tmp280(.YS(n_1798), .YC(n_1799), .A(n_1478), .B(n_1650));
  assign n_1830 = ~(n_53 & n_28 & n_1217);
  assign n_1831 = n_1830;
  MUX2X1 tmp283(.Y(n_1836), .A(n_1728), .B(n_906), .S(n_739));
  assign n_1837 = n_1836;
  HAX1 tmp285(.YS(n_1842), .YC(n_1843), .A(n_1734), .B(n_1729));
  FAX1 tmp286(.YS(n_1848), .YC(n_1849), .A(n_1740), .B(n_1735), .C(n_1601));
  FAX1 tmp287(.YS(n_1856), .YC(n_1857), .A(n_1746), .B(n_1741), .C(n_1607));
  FAX1 tmp288(.YS(n_1862), .YC(n_1863), .A(n_1754), .B(n_1747), .C(n_1613));
  FAX1 tmp289(.YS(n_1868), .YC(n_1869), .A(n_1760), .B(n_1755), .C(n_1619));
  FAX1 tmp290(.YS(n_1874), .YC(n_1875), .A(n_1766), .B(n_1761), .C(n_1627));
  FAX1 tmp291(.YS(n_1880), .YC(n_1881), .A(n_1772), .B(n_1767), .C(n_1633));
  FAX1 tmp292(.YS(n_1888), .YC(n_1889), .A(n_1786), .B(n_1773), .C(n_1639));
  FAX1 tmp293(.YS(n_1894), .YC(n_1895), .A(n_1798), .B(n_1778), .C(n_1645));
  FAX1 tmp294(.YS(n_1900), .YC(n_1901), .A(n_1658), .B(n_1792), .C(n_1651));
  assign n_1906 = n_1670 & n_1659;
  assign n_1912 = n_1670 ^ n_1659;
  assign n_1920 = n_1682 & n_1664;
  assign n_1926 = n_1682 ^ n_1664;
  assign n_1952 = n_225;
  HAX1 tmp300(.YS(n_1958), .YC(n_1959), .A(n_1001), .B(n_1831));
  FAX1 tmp301(.YS(n_1964), .YC(n_1965), .A(n_1842), .B(n_1837), .C(n_1959));
  FAX1 tmp302(.YS(n_1970), .YC(n_1971), .A(n_1848), .B(n_1843), .C(n_1965));
  FAX1 tmp303(.YS(n_1976), .YC(n_1977), .A(n_1856), .B(n_1849), .C(n_1971));
  FAX1 tmp304(.YS(n_1984), .YC(n_1985), .A(n_1862), .B(n_1857), .C(n_1977));
  FAX1 tmp305(.YS(n_1990), .YC(n_1991), .A(n_1868), .B(n_1863), .C(n_1985));
  FAX1 tmp306(.YS(n_1996), .YC(n_1997), .A(n_1874), .B(n_1869), .C(n_1991));
  FAX1 tmp307(.YS(n_2002), .YC(n_2003), .A(n_1880), .B(n_1875), .C(n_1997));
  FAX1 tmp308(.YS(n_2008), .YC(n_2009), .A(n_1888), .B(n_1881), .C(n_2003));
  FAX1 tmp309(.YS(n_2016), .YC(n_2017), .A(n_1894), .B(n_1889), .C(n_2009));
  FAX1 tmp310(.YS(n_2022), .YC(n_2023), .A(n_1900), .B(n_1895), .C(n_2017));
  FAX1 tmp311(.YS(n_2028), .YC(n_2029), .A(n_1912), .B(n_1901), .C(n_2023));
  FAX1 tmp312(.YS(n_2034), .YC(n_2035), .A(n_1926), .B(n_1906), .C(n_2029));
  FAX1 tmp313(.YS(n_2040), .YC(n_2041), .A(n_1676), .B(n_1920), .C(n_2035));
  assign O[0] = n_145;
  assign O[1] = n_78;
  assign O[2] = n_22;
  assign O[3] = n_352;
  assign O[4] = n_1365;
  assign O[5] = n_20;
  assign O[6] = n_415;
  assign O[7] = n_1676;
  assign O[8] = n_1217;
  assign O[9] = n_1952;
  assign O[10] = n_1958;
  assign O[11] = n_1964;
  assign O[12] = n_1970;
  assign O[13] = n_1976;
  assign O[14] = n_1984;
  assign O[15] = n_1990;
  assign O[16] = n_1996;
  assign O[17] = n_2002;
  assign O[18] = n_2008;
  assign O[19] = n_2016;
  assign O[20] = n_2022;
  assign O[21] = n_2028;
  assign O[22] = n_2034;
  assign O[23] = n_2040;
endmodule


// internal reference: cgp-compare17.12.mul12u_pwr_0_709_mae_00_0109

