/***
    * This code is a part of ApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under a XXXX public license.
    * When used, please cite the following article: tbd 
    * This file is pareto optimal sub-set in the pwr and wce parameters
    ***/
    
// ../../../cgp.nn/res/11b_160129\rcam\e10.0\run.00042.txt
module mul11u_pwr_0_159_wce_09_8461(A, B, O);
  input [10:0] A, B;
  output [21:0] O;
  wire [10:0] A, B;
  wire [21:0] O;
  wire sig_25, sig_34, sig_35, sig_45, sig_47, sig_48;
  wire sig_49, sig_50, sig_51, sig_52, sig_53, sig_155;
  wire sig_166, sig_214, sig_215, sig_216, sig_217, sig_222;
  wire sig_243, sig_244, sig_246, sig_247, sig_250, sig_255;
  wire sig_272, sig_275, sig_278, sig_281, sig_285, sig_292;
  wire sig_308, sig_331, sig_340, sig_343, sig_344, sig_354;
  wire sig_359, sig_360, sig_362, sig_363, sig_366, sig_397;
  wire sig_399, sig_400, sig_401, sig_402, sig_403, sig_404;
  wire sig_406, sig_407, sig_409, sig_417, sig_421, sig_424;
  wire sig_457, sig_458, sig_460, sig_461, sig_462, sig_463;
  wire sig_464, sig_465, sig_466, sig_467, sig_468, sig_469;
  wire sig_470, sig_478, sig_479, sig_480, sig_481, sig_515;
  wire sig_516, sig_518, sig_519, sig_520, sig_521, sig_522;
  wire sig_523, sig_524, sig_525, sig_526, sig_527, sig_528;
  wire sig_529, sig_530, sig_531, sig_532, sig_533, sig_541;
  wire sig_542, sig_543, sig_544, sig_573, sig_576, sig_577;
  wire sig_578, sig_579, sig_580, sig_581, sig_582, sig_583;
  wire sig_584, sig_585, sig_586, sig_587, sig_588, sig_589;
  wire sig_590, sig_591, sig_592, sig_593, sig_594, sig_595;
  wire sig_596, sig_603, sig_604, sig_605, sig_606, sig_607;
  wire sig_636, sig_639, sig_640, sig_641, sig_642, sig_644;
  wire sig_645, sig_646, sig_647, sig_650, sig_652, sig_654;
  wire sig_655, sig_656, sig_657;
  assign sig_25 = A[3] & B[0];
  assign sig_34 = A[4] & B[0];
  assign sig_35 = A[2] & B[1];
  assign sig_45 = B[1] & B[8];
  assign sig_47 = B[2] & sig_34;
  assign sig_48 = B[3] ^ sig_45;
  assign sig_49 = B[5] & A[1];
  assign sig_50 = sig_47 & sig_48;
  assign sig_51 = sig_25 ^ sig_35;
  assign sig_52 = B[10] & A[10];
  assign sig_53 = A[5] & B[3];
  assign O[14] = sig_51 | sig_50;
  assign O[10] = sig_52 | sig_53;
  assign O[6] = B[10] & O[10];
  assign O[0] = A[3] & B[2];
  assign O[2] = sig_49 ^ O[0];
  assign sig_155 = A[5] | B[9];
  assign sig_166 = A[7] & B[5];
  assign sig_214 = sig_155 & sig_166;
  assign sig_215 = A[10] & sig_166;
  assign sig_216 = sig_214;
  assign sig_217 = sig_214;
  assign O[11] = sig_215 & sig_216;
  assign sig_222 = A[5] & B[4];
  assign O[9] = B[3] & A[9];
  assign sig_243 = A[10] & sig_222;
  assign sig_244 = B[2] & A[1];
  assign sig_246 = sig_243 ^ sig_244;
  assign sig_247 = A[0] ^ B[9];
  assign sig_250 = sig_247 & sig_246;
  assign sig_255 = B[10] ^ B[2];
  assign sig_272 = sig_217;
  assign sig_275 = sig_272;
  assign sig_278 = B[6] & A[10];
  assign sig_281 = sig_278;
  assign sig_285 = A[7] & B[0];
  assign sig_292 = A[10] & B[7];
  assign O[5] = sig_250 ^ sig_285;
  assign sig_308 = O[5];
  assign O[12] = sig_255 & A[1];
  assign sig_331 = sig_275;
  assign O[7] = sig_331;
  assign sig_340 = sig_281 ^ sig_292;
  assign sig_343 = sig_340;
  assign sig_344 = A[0] & B[7];
  assign O[13] = A[6] & B[4];
  assign sig_354 = A[4] & B[6];
  assign sig_359 = B[4] & A[5];
  assign sig_360 = B[9] & A[8];
  assign sig_362 = sig_359 | sig_360;
  assign sig_363 = sig_308;
  assign sig_366 = sig_363 ^ sig_362;
  assign sig_397 = A[1];
  assign sig_399 = sig_343 | sig_354;
  assign sig_400 = B[7] & sig_397;
  assign sig_401 = A[4] ^ sig_397;
  assign sig_402 = sig_399 ^ sig_400;
  assign sig_403 = sig_344;
  assign sig_404 = B[9] & A[7];
  assign sig_406 = sig_403 ^ sig_402;
  assign sig_407 = sig_404;
  assign sig_409 = A[1] & B[4];
  assign sig_417 = A[6] & B[7];
  assign O[3] = A[10] & B[7];
  assign sig_421 = sig_366 ^ sig_409;
  assign sig_424 = sig_421;
  assign sig_457 = sig_401 & B[6];
  assign sig_458 = A[8] & B[10];
  assign sig_460 = sig_457 | sig_458;
  assign sig_461 = sig_406 ^ sig_417;
  assign sig_462 = A[4] & sig_417;
  assign sig_463 = B[7] & A[5];
  assign sig_464 = sig_461 ^ sig_460;
  assign sig_465 = sig_462 ^ sig_463;
  assign sig_466 = sig_407 ^ O[3];
  assign sig_467 = sig_407 & O[3];
  assign sig_468 = sig_466 & sig_465;
  assign sig_469 = sig_466 ^ sig_465;
  assign sig_470 = sig_467 | sig_468;
  assign sig_478 = A[1] & B[6];
  assign sig_479 = A[8] & B[8];
  assign sig_480 = A[9] & B[8];
  assign sig_481 = A[10] & B[8];
  assign O[8] = sig_424;
  assign sig_515 = A[4] & sig_478;
  assign sig_516 = B[7] & A[8];
  assign sig_518 = sig_515 | sig_516;
  assign sig_519 = sig_464 ^ sig_479;
  assign sig_520 = sig_464 & sig_479;
  assign sig_521 = sig_519 & sig_518;
  assign sig_522 = sig_519 ^ sig_518;
  assign sig_523 = sig_520 | sig_521;
  assign sig_524 = sig_469 ^ sig_480;
  assign sig_525 = sig_469 & sig_480;
  assign sig_526 = sig_524 & sig_523;
  assign sig_527 = sig_524 ^ sig_523;
  assign sig_528 = sig_525 | sig_526;
  assign sig_529 = sig_470 ^ sig_481;
  assign sig_530 = sig_470 & sig_481;
  assign sig_531 = sig_529 & sig_528;
  assign sig_532 = sig_529 ^ sig_528;
  assign sig_533 = sig_530 | sig_531;
  assign sig_541 = A[2] & B[6];
  assign sig_542 = A[8] & B[9];
  assign sig_543 = A[9] & B[9];
  assign sig_544 = A[10] & B[9];
  assign sig_573 = A[9] & B[4];
  assign sig_576 = sig_573;
  assign sig_577 = sig_522 | sig_541;
  assign sig_578 = sig_522 & A[3];
  assign sig_579 = sig_577 & sig_576;
  assign sig_580 = sig_577 ^ sig_576;
  assign sig_581 = sig_578 | sig_579;
  assign sig_582 = sig_527 ^ sig_542;
  assign sig_583 = sig_527 & sig_542;
  assign sig_584 = sig_582 & sig_581;
  assign sig_585 = sig_582 ^ sig_581;
  assign sig_586 = sig_583 ^ sig_584;
  assign sig_587 = sig_532 ^ sig_543;
  assign sig_588 = sig_532 & sig_543;
  assign sig_589 = sig_587 & sig_586;
  assign sig_590 = sig_587 ^ sig_586;
  assign sig_591 = sig_588 | sig_589;
  assign sig_592 = sig_533 ^ sig_544;
  assign sig_593 = sig_533 & sig_544;
  assign sig_594 = sig_592 & sig_591;
  assign sig_595 = sig_592 ^ sig_591;
  assign sig_596 = sig_593 | sig_594;
  assign sig_603 = A[6] & B[10];
  assign sig_604 = A[7] & B[10];
  assign sig_605 = A[8] & B[10];
  assign sig_606 = A[9] & B[10];
  assign sig_607 = A[10] & B[10];
  assign O[1] = sig_580 ^ sig_603;
  assign sig_636 = sig_580 & sig_603;
  assign O[16] = O[1];
  assign sig_639 = sig_636;
  assign sig_640 = sig_585 ^ sig_604;
  assign sig_641 = sig_585 & sig_604;
  assign sig_642 = sig_640 & sig_639;
  assign O[17] = sig_640 ^ sig_639;
  assign sig_644 = sig_641 | sig_642;
  assign sig_645 = sig_590 ^ sig_605;
  assign sig_646 = sig_590 & sig_605;
  assign sig_647 = sig_645 & sig_644;
  assign O[18] = sig_645 ^ sig_644;
  assign O[15] = sig_646 | sig_647;
  assign sig_650 = sig_595 ^ sig_606;
  assign O[4] = sig_595 & sig_606;
  assign sig_652 = sig_650 & O[15];
  assign O[19] = sig_650 ^ O[15];
  assign sig_654 = O[4] | sig_652;
  assign sig_655 = sig_596 ^ sig_607;
  assign sig_656 = sig_596 & sig_607;
  assign sig_657 = sig_655 & sig_654;
  assign O[20] = sig_655 ^ sig_654;
  assign O[21] = sig_656 ^ sig_657;
endmodule


// internal reference: cgp-nn-iccad16.11.mul11u_pwr_0_159_wce_09_8461

